`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IVdnpZhnI44pxLCqFnlTATeEWtKV92//SJ3+lybjGzsD2ofK2ZFkVAZVNDXKgvNdzFz66IGOnVuH
VLHW7u0agA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lcg/Y2fd5bpn1H4GhNQ1sqV0WGQWVmOa2qrr0MJGA9ldZVPHoBiTk++hr+34eTUs/Yy5FtRh/iTb
FWhZoJ+zGJY3eRb1KpdH0NXxuLxfUCAddlzQZmjZygI5w6K+Ntd3FxZlKlFIi8mjVeEcdG7CuSqO
Vq11NQPalLlvVw08loo=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
drA709V5XMsFiNUu6h1fPC5f3kI2TKVu8UDWke2470ztkJrPp+L521NPXDpJJAMj77pPw6iORM5X
RXMEV5QVXyu/Tc8dBSnCzmelYF+n7uuMdYbZUBzhoND5FnbkZPrG1O9athd6VJllR7SR6Q5njjTA
g8NojfvPzey8A7gXAKU=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OZHkbEiLy0CAuNG6gVwPm/NBocxj+JCAkC/cAG1R1Z3osCyuo8QcvaMwmP0aDRcSAM8trrVXNcLx
qFC/Jolm82ryUF3pRO86FiEJYjBUYV10uR7bK8xpAItZjosp4E6Ndi3SkRV3kWQHOPTQZVcLLkiy
rEdCABB6c2sPMpM/6P4DDfgvsz+PkaGIoD+iSMhrR0mKjMFvWvVSuixvokT81pdXtXKu0aWStYTq
BwBSnxrd62iRgRmT8by8XBjs/F++rQxC6oTUPH4RXIiMspkF5+gdMB2CcDRkSqc6UcisYVgepftl
ahY1dPzkgcJx7Rj3tSrNaZTz2kziM8/M0JMcjw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gLf7ExRz6U3DRoiuuOu0DFmAbLZOdOFlVhjaBqXGvtD+RxroAzSEtMsOx+o4fepF8BXkDQKwF7GJ
UQkEZ+zNgGgdn+YUsCXzJ34+6B8CVznOGpblH0pcNG/dLa2An1wESPic39g1k1ak+1c93JW9cANV
plqJ95qtqtXy/CMMAP1h2YS4efruw+gClK34wVLrs3qebX3yF2BB+L6yuaI4IdonaP0E2nTF49lB
0vSnL/Mc1k8NfMy66i74dTrNV0iiLgYcQhQ6I3hjOQYzlcCkvDhsOgj1UWJ+e00hujHe5DQoYyCK
761Nvki7D86KNS4veEcAjjselW2Uu8uSanousA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Xe7khjdGDRG0yPcJxAnWeZyIZhwGiYf3BfUh5EOZoy7Vtgaqu4zE4G97B81XSifQNB0iey3Knvu7
KM2YViDXkptxr2xVU7li1A0fkaiYZO72ahaw5mKUeV3Vkazys4sTcjboIx88/mc9WBPgly/YMZIE
w/bBXuiiUKW3L1W2hn55jUPuMz4ms+r7+kImBkorjY3dtQ+O1FcLwhtx9Aj0NZodRXm0x+2mLIiF
8TjhFyEXsMQ3Wv04MewRvMsigLjuV49fLK3YMtlii+t3QP8DqGUDnnlhGq1XVYvjb7dr3EsIt7+/
gh8th3rL2i4nShsQcV3OPQ3Tu+a0j7ZVr3zGmA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 63104)
`protect data_block
ABT8MfODbmfYGdvYEchk0Dwcv/fgXFWEt3345OAejkK0VSHWxUZMeQMt8f0tBnnYyAJLp1QfkuOE
thD8y1YCAAi9uhksLeEKOCGa620O8jB01NM1qg+fwlXS3vEb03DPb8raSvE/fsJ64vlQznLKVKyF
pMtISL9OSPPcuHanfRrpsseURj4pNxYwrFiytzqn1QkAw+7g7at+JdpiNr+kZUKALa3bg9YRcRAe
e7emye0IHXg/dBRBd0CYgZVQnr/HI1mVq9XJKk02I4DH9djQ+fC5ua60xrDAXmNM83qJlHqlRkUx
e0lsvJoK/hhtVeuqVbTwIlkNdK+lTZkeppyBlxtv48YUH5Apzk9DdoLBPDbv7CNA+4jWUfSEH0N0
RxpKWnXY5g21ICH33VZiG7vN394fvMr6D97iMLOLo5UWbbNrUJP1U2TDJvPw931Cg7AkCWyuVb6h
0XJkQNttFsHZfPmTl7Frsk1Rw3pnuKn2bm6bE07+YYEcbmqHfJya/zJFyoWWhqmKL1orqwPoXzCg
ty5396CNntKFc7NSAXwhVSqsJ3DmjkkMBwAiFhm1eiHnl6zUyosclLB+PWt5zoMg71g9G6lV0HTQ
VYZtcW3igKHDlNYf9/fwtzSn9HdWG4sYdEe3szW4nOfw89aUyh/qoV65H8nMim9sEmQ1qVNH8kw7
28kcrfoFwDVlYzFmzbUKUCqreWnQKQH5Wswq7e0CCEPRR0AOi0iRH0Kxkl4301heD/J12OB8Z4wb
SOgVVH0PbeUSN55A0UoUKNd2dT4AxPkEUQIecWefHb4jF0mQggu8Zey+Nxp/PdelGK1/ulcRjees
N3Xv+tqr3mK9W26vx9aIVWGH2DNl2dyESBWD73B8T1tOKoKyqRtuMnLK6EMBZFSsEkIpMBsTn+vL
uTlFa6wd1bTYGWFTmkShLHr4HaCiTWOOqcBTq17jJxUXIrhgxVYq3SDLoka5cG+RpgOW0r1tc0KY
o9UnmrTKDv32Z3SBtUZatVNtXE52IBIwhfdLXokKN3p9NsxKiVxy/odMV6jCmdR/Ev6xT+qOMC5X
sYw24Br1RD1Wi8dHPjnf+M/lZ8kPOIc2NieKvjLsfXM/rWzG0X1iaREinXVsr++qPq+qs1XxVR8J
iZk6ySB6rVw30ZX8PlxInX/0PMm9JpzF7MD8fowHKen2tU+qGQ/CVJUaUIgn5HA/5iRL6b2uOR1G
Jb+T+A6F21h93EvjL4spSxflsZIEKnpR9mXOwQzwADldnDFJpUIuM/knps0DQwxQMOM17jBZSduf
SJG8N5f7aA+3bxa53/QJMhBdK/K1J/j6n4Z/E2qvdbhbw0ysdihqlBnsnlmJMZZnJLn5pVYvkylN
szm+3zhAd5o9Q90FzOoraLJMUDYmmJwCCYDclOBa3B1I4KDzBIFwC+vkPpQunyzC29OGVovbOnId
ltyriOgnZIbElP5EM/+fEw3v/GU8dd00rgLSISZPmu7wVWptoeQz1ib150Am29v1Nj+O52oUIp5X
c/qGv/vjZ5yphknl81rwGB7bEU/YAe51ChiDArYiJ/Zsb4jmM5HtLEimRNegpTFM3C0l69iBEAnX
0d67J0UUfrhMAHhvgjyS2Tabf7kaxPQNnBrJ7SjWP1Zai6HviazVb2j69YFDJe6g/E/1LtZNzCl2
TXOgIgYTRK7+aIUITfOJth4wnfLyuFhNoqdCCZxkB/xlWP2gawTIhMvO8U+eHnIRgkcRJ69RcHlS
wUwuve/m6PJiHLP0pHjOkCQmrvZoL2V2b3+j5k/UCfFd0cpZ44U3Iba4l6KEoyw2rHnfLapl96Uw
8tpBgEm5YEuo5xL6wTTy1qNMkSInODv+i9V6WS46lBd/pK24r/nW8ExbY+E+jn8b/tDIJCelnQX/
g0OeLCNUXOLP5ET5vha8z9FfMqMKkjDs0QgAfNhSnt+2RqLk2kAPfEU1pxZV2Bj3OIyC+QrHOOHd
xTb4w0lcJ0yDkT+anHuxq4TeJDFFLWsnpaC/CWEPMq7tw3voeGCccWNQIHrbyLSq2iFjY8cnne5o
kalyI70YuY06BLd4vfF+JWa4E9ZUsngfioyic6XsfsWj96cpTezjd0cO3mn0wFuMmgXZXSJo1cGg
YdMjYTPsHVe2aoCr2GZTyfGTgdTTYjWN5Xow6GqG4ltvSH/j0kCenOKmhnc1QVxwX1O/x2Gb/MUq
3Z7xxSnBdEQmo9xXrz6ruagPi721+Ru79xSiXiVl+SKLgeYNV/1DXOm5srfAdVQkmDPVjpvkg+QS
ofLSrkiT6qORHsf4cVuihpN1BTt256HbsU/UXOr9M3BsyDoc8RpjHDCmkoRf85r5p0sQ96nIjttr
3tCqQHzvyMswZBZCAaL9ZK+cA/T5V7+bA8XRxjvl+QdW2RIv2PeNEbW5MbxG6hW9VVl3dP8GvqtR
J6DmNfH+QIAXo/kIs1zeu4w81qmHSacul4741CSUm1RipaKems7aSA4fwPnaMGyc5DWYz8t0z+2H
HgvV4uOy+Rd0F5UMKmOv8SgvhI7P4jMHQhMmhWFGl5fYQlBWqqembLpj8AczhxvQtd7Yauz2Nl+H
XT84jGfxXejKinSb2Ah0FQNxxd04MuyqgCQUJ0cT8EJykgZ/yD0f7AcQXaQ4W415CfmA31OcbWrk
ZbVAEtTZxMgzaqL6hlxYCiQi32rzs93x3V7d1pCnAB5jnCOlZjZYwmcPVTVx95RulqRtcamrI7QE
zG9nmhs+JpxDCdUKQH7UkDq3keW8k8Q/qVARa4BwqdIQA6fl8Qvzcwi4+OperCVjiNd/rCDbrlxF
NwNGgYC+LAFVDQJRKKo6pLWuZwB9iRb7s8RmjphcsJ6pjf6H/VO8hGb3z6N+Y+9iZ5wjee8KXzjz
yYIYNRSTJ0498xzzovgRMLFct3gwxf1WJpmCpnXNFqpBcGGOpc/484wrXhN9IYchUCUx3w8Q0mRJ
Kn9YtDTukc8+5M/yJXQ6tIa2nI+Oic5i1ZrraY/1PCIi3dJCVp01hrL5CdCJ6us0eI5wbT7A6JXK
G1GO5eLshIBTByMmHUJOfQsD37h0kVJU74/ZN8QqHSTCZGZ+eJd3dBTKEl/lvQhDIHqzRVRn+QY0
HtQkuZKyENcI0chjZgyV5cQ7mY8sNwDZvp5rjoAfeloa8OkYonl731RlqxzvQBZ7/q+ca38+lta5
EHMYsjnzcQP8XeO5WmHTirSS/yh+tZWfRnkGDGM4Xpa0EbZwvardPw5DF63f47hjuAYuq9EY63ut
oT6vktdRmLBuNw/t+xgf7lOthS/dk8l1/aPrgXhTYwWFFkN8/OzqZs9IJPg71PvRVn0yLonAyMVG
FBvQbEQK1eJQ/Z1iD7MpiotiVNRExj0ycqknrSJOGCKmCCTeBf8MoV7iNi6DEdSkw6/NSIxOpngN
IxB5VviXW2SNXZ3yVoWX05bdaMyRR9SUsXvQ7tAbET7NAt/6k7oJK7LeDW65ytumFnjrpC102Hd7
zJjgsrjm4zPL+ta8/LRoNAbm4gF2HVx1GR0qJ/BlmA3sZfzEXVcf5+9X4G7k2xGQa42ijVYqIVVc
iJTY1K9HCq/4FxHvH9K/nAgiMZaXgv9wxXmYF6UzFa+RpfHvzM86eRjB4H9yq2ITM6ZlN4MEBcBI
Zy3uIKAosbGcpsF6Zbce+QgS1HASczbEE0M0epYAN2X6amSI7mujO4C4nRlE3w3OmdD6QRFG8AwZ
rF8n+QfFEKKaG13K+8iHtfGzQT2KEo+WjZjRJ8YefQLtvORr7lzyyl8uYela5DAA+h/Qex9VVaaR
f1KD+NJ4fWYf4rYrGvSE9xYUgpsNTvOPMPjAUJSwa+bDPipRSwwOlo/x2p6VqVl5cE+q8fMx0+Au
9qY65HKCx6VrBsqPvnk8dJnP2X1JRtUp315ZGFVf8juLAcgdR5Mod54w6L3LU56To4G+lfP4u1Pv
kOIdqtSeEYAh90LpIc700WypMlORibrkV1KxPtpKAr+HXA3P9IV0heWdvJ8DvNdJxLXs2utO0urn
JXU/4K4BKfxRdTM255nn1dChio9MMYpI7wG2ZYdrcZdeLoABSWx401jgg5JnLXaHnHfrfu+FtyMw
62mmIHraZKDrsDuRKtlSHuFunV4cbRcNc8fCq06m1gJE9+UN6devlf3QaMqup5WProNmvmpIdirO
vZszfAEHInTD3msU2g6DfPFlP1VtFTn1cwKGd/vCjahuCLYxA01y7OT2FfqkH5Wyg7+yJ+NtGMte
NW0LZllYQ5OVkifeOvisONSrt6JO8FYsp/XUF4yLXCEDdS/ub+lSM5oat9T5LDRCg7PoZlbK3S9r
yOcLyulAahM5voNJTemtsANFqlGEXcAsomZMx6VwPYiO06dLBJWC3RyCfU0ZKR3fNAdDJWJDdKW9
f9xBApf+kFKFHUu2XvsxH3sFAodMD8g8EUTzOgx2Rb4W2fHz+Dpxnt2tGZiSiQqVzk1LT5Clqd4j
nM4hQX9/P5h8h1Ia9nACm9uZTCkwjz0MLAVufBQw2Hq53ZJPrJHTpJPbehkd8bhrT3P9nJIw6XcT
E8yaHynaIKWzLxvsytluv4SX6V+jf+4NGKlvi8WRMYLvTu+D+NBQ2MqQTBcj8AcPiQfPnJt/C6t2
+sLzLZIU9I/78D5oDlJXbd5p0fljI6PCPFxkBBIStK0mFHkhUNWUgZ+EN9hehNrG2dx6kh0jzOMX
YraE2ewQRDxMLxUyKLF2cciET87ISCinqkkdx6X7PEq3mZCy7nNWgVuBxhsafaHkfy1VLn7sehau
T7taPCpNDDZJ6rqc3yNgXjqicNikwjDbxGTE7NdSnSTKI56LXMxor8fkRxATxDuZ5CD5x+Y+1pzi
QO4A9Tb6myPNiS+OYPaIePzLNhCH0FpnFkxl9wrbbq4iPwibbA/HbEatMZ+IVtewv0r64m2vq+HL
jb/xgWhxGRIoE1/RWXvbJFiuWF0Ph6zPVgvqxz61xJojrJtPsesU8ytNwNNVULoBpqRVai2L9HVq
NZxczyNurt+JVa+yhmBie9Mbud8P8YS56RDHnNUd2ZA+W5UKxCfLVtUCpp2nIUnTzIbk7K7Dncnn
D2L8pFw+q8Jrn6U5XL61vszDZiPidnkIFEIMSkVzVGgOb4akGkN0WqV5G7LrRQdbHTWIGBA3jn5+
OU47a2LHkmVq37pNn8uHfKsa+nnZiZzzAZHzfOfSAc33CeppV85sIaVSVK8fjYMusEuE0Fq/i4Nd
APeWUxvMYxYqFlkb8W/Szc4bbjM720UQ4g1IPj5k/sudq5ugJh51x5ee1umOuIc9mSVqoBs63I5z
xJ1ZDKhutootmPXgKb/HSU7Nzxv/tj6BAnmKLZUGe1wBiTbKHgVc7R86352dStLA5MJWJgvVUR+a
Mlq7dqwxPSdsnw/eh59JsRNYp+mgUTeZmAtqMdubE0nvK7Z1gylmXHOKjZKW+vmXABQJJaga8btz
SqV+ComZcoPy1HaKEPhAisdE5EX/EFul6/SKWetjv+wmprekRZwxfxF9Lymqvf2B7wAuaePPmwRL
LqfpfFwMP0k4bagMbFKM5+GPA85YmD8DNN/KbjCeEMLTYpTBvUE752p2jAeIP2YcA23srqmdPKjg
Wqsdk16N0Pew6TiJ6Q/KEptIXYhXumqglZqn3YxUOj/Cqrt4r0cIAsczTzt+9DwpjvNY/ruAhfW2
AIS0XAw02pay1+1M3EHFyzPUuDTBihAYgPY+qMwJLzTPV2hXkZXmHfXgfHeZfY4CG/AQLy1Y7yOw
VYLv6lVdCHfii5ct04M7vvVMkaBJ0gyA3SaZgYVYZG86Sz9bd7iZJvFou98/8h9fUKGYpKZcrHrN
2khl1BxnLdyF5Qw4Mm+T+GeBB6U3fjuv4NdpGVAbQ7rEFX2dA8Hy8nIkyndToeLL7Xia7eTI2N7C
FzGZYIh5JGAPJiqg2/Sq36N37cffyoTGAV5Yi/mOxt88o1BxfhqFmxTtJTBw2eIqILPAEYKWmtwg
Rof4sHZFyGATHxC78NAaWcHPPtdN8UWEBt6OqrRKohFC5/KXgzmFO0XsCSm4yeYmKxE+gmLmRaMD
SZuqneehvqVbe+vEOlIA8Ss2PE6vPHPuwTREL/RqqXToeepXGdgGyWufV1Y7eAz+iPlKW6E8aGwA
HK8J327s0esZseCNGAxKaiRe+JXBGkclZ0xLajIDpvv21bttxpzimCqPrnoYFvQ5ClMmYgPbyYR2
krRL6k8DL5WkKOafMVhVh0jdBattH5H6cfpbNkjW32GyCaMlsmwWvx1XKmpaI854GSjtW6VmWsvX
wBAZpKrj2bYR+NhDhtUwIqaKexsMmvO6+CHQuOh6tD1y68hkKhUGJF/HWfVcm0EunIHPCPOPJvyn
ikmEb5g3Ijb+9WKR7UlkwAfhegZlZTYSBf63Tyrrln5DR+h2Ie0OvHTrc7kAnpldXbQS0g+JsNjh
BNyHkZXwCeMDx8UKmAfYN/zHf/NJWROBSbImy5J0ooRaTghIlhMbWKbvWGM4Otm3xJjv0aZ8UhBX
0L2tZh+lZSri/4MhF/XEc7DywwJ+3E88d3/IedrmrZvy0qYqT5IU0kOxDVGGfZJqw8pJFQt5XaSj
OQjzbm+Bf/j7Kl63RdIRwtscgqXHGkuhv0LDzECPLFL7qalrs/g7p3SAl/K6wRKBYqqj4gKHUKG5
L+yUKJ2w5UgBEuVsKDc627fTAbCN/qCXUGJ+yI4nhspQW9Hw4ReJAhq08DqtbN/IgbX+YZbVXNyg
OgexiXaF8T1y0jX5n3WrzhW8MTtHUPxWtCr0EQumKG4mjRJR2zE6TI/JIKKy1In7/RU0QiQ/xwk7
ipXtZ9qNexX/ngPf2wDKgAndK3U5LHq/cnESweGQa3DEkAaCYW/pMJWdo8RHj+lHyCx3wdj06Kd8
euerCtgsTWUykeKB84FixqYJ3f30CqRoH3JJLs1YNJv1RwDZVbFXKOEe7N8vKMBdUyQQcLEsNzQP
9uGoV8EvpeFfvjsGfvU4Agod8hsqeTFw3LOFTGAazt3byQZvx6uSCX0y4xc1FMbVPKnHnoZuEmRw
NREvnM+5Vs3yJMjMEfhCxKUVEM1IZtwHCFx6DH8vOGyLLgyxkbQibzgTiGlftIEzIvkiyG6Qhtdj
2qOJiv8btTaoHsYFq3UMUv0O1i2GvgF3WDfii+1v3BhONTAmrYC2qajH0Km8k7BHmMHlb4diGkZr
byZVxr5TFNFwRYk1TdZQGzQj51+WFS2ukCwcEQqYiKwp167g0Jo0hRWAPi2U1iJXS2JT1rTDuI5Q
uQbLQa715xPinR9FEi3wSRsxYW3iU8HyuR5+rIIiVaLYgbvSHWNhPcIREOayozqDIuUPC56VNOSw
4Lfq4HmZU85e7bXrvfNn24+gMvi0FjlmjLq9/xOyLL/Y3WIxDW5o0ldZAOcOlvjTYdsghMAY6YOI
sXX+mLbWmpLuGhSbEI559YU1UiS7IffUlKLskF7tSoIfCWJlFhUfJ9qMltll7ocDI5d7eaOe1ix4
tfC2ekzYXTv0NmLSimYeTYEIVr4M5t2Trto6EiOyWFphlX3uetv1ymvl9NMK9KtJf4U/bnTW00mh
R1EtbV/sQigWs4gubr3hcn4TMW706nu8b3BGMt/l65CKvmNi0BOnF2OheU3r8htIN9dowF+HtdLG
WQbhsvrf/vE/CNJrpTYYfKFplclbf/1mqGsKT01xXTZB7WG28kFaSKCp62wGzK2hf57qWiXvLEaY
Pc+TS6ynSdVv917Ca8YZFF7ACk0L0SMqwzUN5BLDHpgyHHP5Oaei7agw5MRRLcThX3nSvAg8NZvX
9qhqXTnfAap1r2loE7tyiDRVtRvnoJmbCvNDMxL2C10iHCC9tNo4oCLIqp7pUwTqXVZwnMWJolG7
RCphZ8rlJ66+IkwYHHb2St7GLBHarMt9Tb44H8ml+8iQ+dF/F4dHadKXl+TzCKsKZ7E9vCRXQXGs
V3TFYqcSRtobPNDITmTMraTYxo4o9cB1l4mB/dNM1Xi49x54yG/Zv92Mnq/R8beCC0xIpXBxaxFi
PZ9ZSc2oTAEtaaN0L+3sXryldwCtH+or6lJrchUsnpR2o+5OfwFxSyaULCusBMtPweBLyfNVQK5G
ci5bGBPLIifOQhFRXCwYV+Oig+9QUkl4VhnhmMST4qyU6gASCJdXP7EzkoR6/pNtP/Bd95lLGFhF
K18RQm7zcIiXeEQDj+xp7b6X/u5Ut9r8sYbJqRiTLPuvQ4d9KyzOiMJ/dK6MZoM8gitTiO2yEPuY
PrdQL2RrrpajP845Y+1Qyu/JZkiVQ3dX4qOVE/Neu6kVMwqrkJNn4pCigeIT6oOZcPbdpuiQ5mfB
nIy35GhZIbDrZRxKSQipe7+s/1CVQLqXc2B28VBqD9Lk6tH0MXHSUCd1U0/fHXqLMMQWaAmilY8I
/CxCdQ1N25zcdau6WMVKUkXH+dBrWJ268qrtstpbiw7yCH6f3vkTUUyGtGgkEFJ6dRze4jtIW1yo
pzTaz0SADP17fKCJgkazuS7XO6OE1U8OyHo0GIIw+uVWfpPqxh+IZ6MJoHIZLanwfItgTgwZRSS/
G5Ld5SA9h1gChPp+bXaQmVMWOQ33xhwYWJ1HsOqiuDGnNC3Oj5QjNBefIyWNKWaHN2umpncW1xJL
R5i84P5OsDmeTwv74gsFMyFw5qC8Q0l/6Bc7BJS+g8r2P1mYwTwZPDyYbqKK7yUvXQ2iNRuWV4zo
EebjotZaUvrf0gw0c2h/Lb1DhIRgl+wICAhW7gDvWa3skcGmf0TaizVXr+VnGsN72i1AjL3oP9yn
BoefDkDUIab7CnEbhz//mkdU0YKTh5Fpgqum9P++BKUlCFLCVFJtmN7f3O6tJXvCY67bAJLBvyXh
uBmSGOLWVmxUr4LOAzOCgDUOXJJRYcJ/Q6YwzPh4PQwBc15gM3sG8D82wiP6zvJJyrlzrFmj1bUV
HPafYCT+rnetKNHlbs9qB7ctrcKgWBfbwTb0xyf5RzXAM3ywxZNRrT9Pm8xpADXJrRYn3aawJwwX
eQczRL1DXj29mizdbaFKoAZx2e82zhe5FGeh0xmqmcvPaLgA7ORGk7ml4I6hJ78FXs7MJW5EXUYk
pXoBeG83RkLMUMXSnooUfeNaGGRKVqj+l1aOXLmOtDfU8V3MpxAJMTxD0KVXEplcQJcdsNfkU/xk
CB8WRXqD9NNZaeDbJE9887YynsoVYv16erigAmLQIN1VmOFuuF5h53mnA2qEstpqTUIL5lVV7bpR
9mL4S1r+57yEkh+QDpuyRs6g9rr0jZrgD7eXLvARuQ1lQBhDX1XJEaxrtSAabHqaP0Eu6h9fU5+e
+imeEaF2ikXCfBz8LoBnZx/GsNAccXOxwyt4lxrJpQq69rP9C8zX7/Rkohzv62+7NrkvucZ+ykqD
mMqn8D2fr41vuZ9Nsq0PZlxb7kdfTT11/efUIcRtSL07x6V1eShBJrwHN8EXXCt2672QYioaafbl
W/0RhizFmKjq7P3/Z4BPu2nPs49n5QNCdnSP/Do2BXPc2pHvWQbKbne/jN2qn+2MtPEcv4mkhk3l
XQ25u9sRjgPTFOJSRZ1BPrZVTVu2UF03zqQmXzMrxwyVnno4LGKlrBo002QDeiJWEJZ0h5sdvoRF
MwLhXME2rQOlIFPyucN36RcCIYtmCDexXzkfR5s94YaWRKjzdp+USMIu4VvsviZQWuZdvFLa1bKS
X/8/CL5mUhKG9rsHeqtzcx/ZnGJt7X6c0YZXnP5t0WKS9R0+0+RtHwRb5PXxNsVms6jDY7NUGulJ
5y+qq0mg3Q7SZXUDdeIYRabCGyq0ZIk22bIAYEvDyhO11ZHxjMAo/dLCwoK5AfO70l4ke8/kqgDp
oImmKQHleYQiJs3Wv47hYgH1UaLLG74IHfbvyglzuQvjLV7LiHq8GdiE7SX+URagGMGz/2iBKriH
rO08lbft4B6+v+mwnPbQWjdh2ELoNm+xBbmZxawQD+q6UHJ9Vbys1CiAGD8Qwfv9PwqUUliBcFSu
1Xtjs5rp/kelZgaU1OEA/FSN4MXuhUNWxEVutVDRsaHir2ly+rV5yAIvsGPorbrEhYHH2Ewx2dcx
PUv38UI9erdQnP5SrrXqQdp+kLjONLGqMf8Pgzp/fahCUqih6eIS3xmtsJFNxiYXYGhgAnjUzvtB
JIgljyAjqvvihN86ewCHAqYbyA/eQg1uRBoKcFdVyZyZRT2qdXj6SrRgNTAy0Eg5ZjAheGH9obU8
rJR6Cxv/U1KdEPB6++4H4Xpqh8pZb7vlYUlpI8OmTZFVp9yyC3k3u4WFhDw8wSLq9mvy20nOtPVl
pmv5Pz8KGIVwrNTDO+nqZqowcmvNXwNafWCg55HfvELIriAz2pVit2jwqPT69NNfjiMe2ccEjRHM
rAQoDmb2fyGrIgWZHfsJIsOCr5OE7pJLJFOZAYV5+Odvm8PIFt+TykUBkGz6X+oMP1ECsrdyIAtO
o6ryxE93bFF3pm19eFIXbiadzfwlH8BdwytxWKjeqSkzKsch08pcZR0PAHWjO+pa52ucc+whbzhF
5CfeYtNCYqomfq6zK50ZIIcMfrKBusPykes0y7WWmytG7bD4ndxe3smE519fM+XcX+o+kkU2oKNh
18JS+90k2SO47k7GtSSlF6a9+aJm5EbNrcM15QKjylWjrzJ58Alr4OHowvy1QYSLkaMC9ocxe4hq
ZzJ0t5csSDcmxuZzqa3coe8T386ryxEUP9XQjEXYGhxhL8l+97h4ZHG2ZW58ee+55Ws2xlSy/7gO
Q/wAjpI/LhUObJUzXfDNOP8oI2L7cg8xQcQ5S2igBh065Re4p40F2UipHJWv4/nwMLtL77tnAHJy
hyeCgTBqYVvRZa/vrp+OcdL7amwCPuAVMahm9C9JXsHe3+7h41a3hop1Ra77yl4tt9kGd5D1zzcb
u7fbE0Ix9Mq7HzhJbpszff7AQ+9AFBF6x0Oxl+Y+G68JtWT/O/S4dSXKzB4NAPtfxHmFhEjx10+s
AryyJ2obMlZuuo8SNIlTyLUNssTbWptNY93A5MotBoBnqBmeZZv12HTYXyYmIo7XL4kjP3EJs8iz
cgioeA5Y01LSyXYkDrPQXYZWedUNLT2JOzUzDHBcAOQRwYK0DLpzHJIp/Pf3+abfxOmFn6XHqcjc
QElNv9+mP/gDFCJKOTbcgeQuAAgNX8lloP2yc6NV6BXhULkDdXnE/UTmm/Bo7MZxxT/a3ksYphy0
nBbvZqn6DF2izr1w7YDmsyML/gUwreZ90E6PXutGPvHTK0pW6SzbdcBGUO4Jo3BSX2Lq3xJVXBxz
fg4lH0kD726RLRwLezJjNV7XmmAKwR+Kw5+QhBtS4WtKbuWm1tt5pWPAxLtdJ2U9W5YpdpGpe3qd
4agy6cQCUdXXEcx9S3oB9+y6PIISReWtBWE44VSe6XGTATw7N5sUsJtKDOO4JmgSdK9iW8hK0O/k
nTV15j+eSmJGmmTwP6FDQpBNlPyPfKvywsfTiZRC3f312ndzze2weF2bj7QtTDsdipFPPcwOljG1
iAHlSM5rfgfChlmPPS75G2JCTMVpWwzGvNh3rtNEOpLC76JrUkK2CDTG1Lc4sbtfAiqgaucoPpoQ
gUSHLkm9XJNlkVmsvrpdYuTzyuH2mP+mgsCcMteXCplaVySUDtSvIm5bxyK+V3BFE4fznK28qElr
cj37bm6HeDDnY5dYs4dsyn+eKz0SIqQtcWYWByT7vcBJbHuMmaz2eMbe1em3YP/ZPpSdi8aJSyxz
K+UCSQmoz6NtVKWFg5a4CDVnafDnsp8MEbnS5/nVyPVu9otGREAr+x9iVvvJIWjj4fPpoEoCUgBE
d1XeB3+pB2RgEAr/TWTG/MX9/k9RmEQWzlORqhpmLnh3GHxjiMOVh5gBWzqcwBPAeIAQ4Ar7FcZ+
zwo5zrbpvFyRsoV+dudJtlCn6IKeMtqv9Kjyqet5+Af1FlK9hmwi3RuF04T0B3EYgVUwnmPA8Kut
qwn5m3TrN6IaKXrflfdnKQ7vXhYVKmGpttC6jWJ09c/3YM3Okt7DuQB5RmIMTEtcBWsODPaHCPwQ
NmITcQZ/2ZRJ2URISfH4cL7uWS4UF1fPoM6iqR2hfnxcIuiJAGp2ORaRUds4C+GlRDlItoriDIye
RbzwxoThPNKWumCBTyvbDpiTaRQiUcCzSozJwNU4TqsLg5/3UL/0In4GDy3zSHvd/gN5gKfLYBDU
b8GLBM2xsvTkXFuO4ap1ljmOf7RLuKR61VRlsouUca4vLRVZXaqQqy9qwuiYsOaDYCW14WeKBa0t
upIC1mT25zcd7C5gqYq8SDoQ+vK9+C02aeCvRkof5mYz1AEGVOo/1aaqKenszmCq/LJ8y0RwCq2f
475EYvBbe+nl9hLWpSFKUk+gVAeFU34pb1aCnCnh3QAfeimuguK4mEJhmlkhm5k/h1Qz2l7b0+D4
GTb2SL0TaNq7y/Gdn0W11bigsdmgUQ0KI75JkdPR4hJPZzJ9iqXKT96+ZTNuBDXKEiKcOs1H1MFM
zgjs9jXLhtCbGV50E9XnSoerrVU7v1Ehzf9N3/QPPkuHArHbQZtVKrWa/o2zc15ybevZDG+zdSpK
topjhQVgFsDJnA1qfWSRwB3jRwlNSUvCsSQG12S5Vy4KFfiqLXOydLs0p/exvN3QUEkJo3mNIsH7
DA0ianrU10wI1sWX6Jg3JxVhrWSeSbPXgHSvfGLtFZcCc/c0VzdIcz3xYoBJ3ug9fwBDHcYcy5d4
ozfzUaaVVXA5OkL5g8kgt6UuO8dTTETD7N4qZaDEbZtCTlrXp7EtXicCoWD6iTXnOR7DjNWqqd0D
3/3LCoiD8fO3kIqQoWN9rf/r2hVx5FyOWU6I+2ZYxPTUHqTI7CyM4II+DEiRWRHcrjz+Tf8E3Qls
cE2CGXx0BRXMYjXb1V1+9NSnMCMn201kZYxUsf0P9lnGp29dPT0sF1ZvkHyNb6deKO7fR0FpNNsv
zf8kfjH+b0MxlEP7FGdkS4yjYAhM4zugfgGGPIF2Rt3fAXB8PHfPpBputbznTHY0aiEWWMXk6PNt
Y/+FzN/eH6sNsia9KEFqsQ1wfEDZsRTC5A5FPxvGeLFNPgHc57jZVdRZiN98Sj72gYMy9gea5dxt
S9sjYa6tUuABBhKjFtJg+VuP4wmGArC9eDd2voARjN0rv2Qo1ijz9JWUq7k5R1C+GxOvxbak54zA
0RiI2GAXjBTXBX0nyOQujRs4QgU4jWV4/NHBGKY+c4KqVd21WA87yeXVf+mpvKoLx/9NI79gla+Y
/Kt0w1tCaf9JwLAmdSdHjT/yeM7ndiT9yuYgzY4QKoPnvFU2dXk112TLQyr9h76Ts89Nz6Vrglvs
LVSkcLskHPc6YO6Czhw4YuoP8aL8EkX1FucOi28V60iJgZdBEqv+LUaZJM7sfcaM5oPdB9IyohFt
5qA2v/vmTS9s0AwOWGZeihWDzZNgK8QKCrGIKt2bwDAbNYOqzncf0tfnSuaBrTKai8y+WBIqyMFh
E9p9dPvo1SdfDJMq+//v6wZauvrExoOYDYOEAuwaQfq9Ft3oN/5GXp7aqRUYguAqLE3gm2S/EtUd
GIrIdqZcaiadrOKWgn+wJLi/w5ZQ5iyvkPVT8PX0EbM75FmiG7TUR5eG6PSsGf0KLmFWgX/NjFQ+
H0niKya/U/o/9X64AAF0SIY5rzCdgRadfG5pUYtIrt6ZOwfiXgFfVYh+OCWNGdOHPxO25DZMywcQ
0sq761sHXNB++XUOyXX62ieVLmg+NjRQtY6lK5Q2oplx2Tzd3Jpc7S8X47eHM0w20mC6bC3gA4FZ
Z9QqbWcH0kwU+ECkt+quycG/NNBH0+miEUFMKCjnZ7qxVYrkAjTR5ryDxX1DJxb/ioidANlkelcQ
8SCuoZrb/u89dtW0jLyVybBBOcyVPi1G2bTNs2QmNsuaTWgxmf2nI4Tc4zU6/YLoA5tjSpN6ie/j
TenahFH8T+6rXb/UZgY1osXj5QwKQSDtwmM2KwLcNAjxoVJ1GXmcAC+DK7yPneRmnW+vF8/mCfPz
OTk0rcLUhO8SbwhALwk0N7tC6I/uvaew1VwXcDOEQs1gHh71+HZik1RMgCm01PbFarYBe8PZ/zny
ygBWIbnSmkbHnwQBcy3LXnNx7GuZ3V+7CVbqNWpPmpuLG8nnuvzxUVaWbxTiwy1FXUMzzoXAgl55
e1JnP4RSHBg9hQuqla6IsLanZK+6cpIwe4Y17SqIedYTktJzqf88Y368DZgJ8FSE05dRVu3itHnA
mkYXLeWDaB5PpGiGhWOgRPPAq4vv6TC54kLK7pWVBEfN7EMfvqpnWP0r/ida41tXQidOKqvb+TuO
3a1ZxjQMqs4HdclGlpRanES4BJqmIwmd+yiLvoGFWnSJLq5hHwEUKGFEE/xvqzYqCrQgKIOk1RxQ
HdiVSE0l4Cj/X6UjKGF11C96W7UipSlB5oOjTkbTNzm8tioEmmOn6hXBE7tTgrpTGKl3sk+Kr5S/
jaQQ72ek51ctIWArXLQgpLl3EdGoKcTIBXUZS4tmSqFElAeWX3RyRJQ9+AKtpurIavK+gRM5koZb
9YQgv3/W3kwlq0dllDgGIrPGxBZmfjEKwhfOgPAQn02o8oVLbLal9PtSElF7+nIkmv2jVMzIMu36
ERFzP32qwc7GpegAE0pQkCuyfN1U5QRW3DLdv7hz6GnN6t2ssbBxemnjESh1xgOLd1+eFKFsT1Pq
HOVERFcnXPsARSddMRTzQ+tVd7pWC7FKF5TrBZQW4v/+HCA9bbiTVgfcTlR4eQYVMll2QTxaEFDU
xSsFwX8Y3b4UQxKkYGiD90eCpMmUzsh/I8ZVv2B7q9nFB22aZVrmFKlmAMhD9ILjODw/euGLWxe5
sX9xTxLlPKYQ/mTH1zucVSJbHeFMKOT1nP/12BXMCsOPTfRVpQ/FnPTYK0du6mthC4//4Ui/rwKU
JCQUrpUZqkEsKug9w+beArq5hfV+7qpZ/UIyXTvzCnj3SGxOg8a/TqgtF33ApXs/ogJT0A1qTV1u
DXzO24vH70Seeblbr8fTBDBFDtx/LUvXOTTbtQ+6bRYjHZxbjugjZVKrYfzOz2i7rJ+PEXQqELsA
e6c7vtWPyL7egQU0j+pWTJFBWuNeraD7IY2/mNhMlm4uQ/tj6wCtMj/G0FbUPpb83yU0aMI7FnHJ
Vg5oFaXpDCxtX01eu+wcNqQ3Kpy/AXbBfLfmFwIwxcqa0Jw2GxIcU3a0TAiWGTlUUxKLTc5Ihw6q
Z4QB8eLnSowyYTVCfOudu61CRJTQGNpM/mhyUSObPG1s4oBzMuXm4+Wb5yRXPKCdGBvm80kFy840
ig44F/p6NjS2ar0VDQYAIrCQ0+cro1cLdq+VyrIHZVx8WwxK83jbPy2EN4ptAzMkWBbNViXGhS/+
b0C5bKz11MpHSzkDPK7F7K/izFHFTjeFO5baRO2JUx3vwo42Zzj1RVdYo5GugKfmDlOYMe6BUIF1
i0RmWfGylF1aEi8Yc0UZLJNdqzsmIrfNyEXrYSLI7RgxpSf4ON1/gjwRLZehE9vqq3DoO/eEziZe
GsjiLndP3JzG3RHcOrJOM7a3hFx4gVgDrKMtaggAfQqZzMrlrHWCVDE4kz1BlVAqRs4dy5lUj/TX
Pa7FPxingf502OSD9tsGxPku53eOvnqYXvmOHx3tRpv1SRtn6k7S7QhUivg1KlUlIw0eIQyY+HRI
Wy9MfaZHpHuJOa3XeRG732/e1FAKy26PvBsd7sYbYN4t+LbDY7bNBeTaq0oKSUmDnW7CEguQxmm8
SA2UfxIf8Lvz/KbrKFs7ObgExA35veDvlO6lv8MPbTOeFxKcuW6MAo2eXkSzvqY1WxtoOlAD2GEd
P2IZOxzoShDF9WbZ9LiHiRsn2/gb1GSEUkz6usqN3lGPumVsTd93zslrPGUrqTMcKtFcxaet4Q6N
RP4Fe3Himz77SrchDaSBDSBVAA0E46ifPYp69eRoLoogQdRIiHCx3mNDgGySEU+JaM5RZEi3kBey
gu05LCRTtbj6AyTjX+jqdyv1zlqEH9xTHCt/XJHopmyqbETNDa6PZdKR755uTvSHm1gpXnZu9oea
pqCUs4b+IPybEPl/Cd8PnaObvkXQuaT0wxOUEnsTSBX42wNOYggpRpDwG5B01o1FUgcmX0T29qi7
3qZF6N9TTnnNLOMitgv7XwRgoaxd5TKcf2FtoCEHw/HwfdgYTWgO+UbWck/0faqJLUhJuhVlnJ9R
pqBscPDIO6UFA2MAnq7n2KEaP4bLEQiVmaHluAt5IZZCHIwvnbPRhJccg13Zvh9VAo4rJAemEtPE
MTmuI1vKqP5hEQh+NxV63KmJ6lOrQEwL6VjdCOEluuVJFb5l3GZ/jbeXRgEBefSfN5XqpxjLSxgZ
23UvXNh3mKwFzxbjWztO7Uqm8AJg7ZOqG+XMRCOXQVjSUQjD+bpZGfmRnlaWg3wxBVksez5xAImd
EW364tsbnfM1NkQUBqew6MUZcYk8KGTu3pJQLDH8QsLYNSsgL1rh547+fudlRI7J8qmn+hF0qmjP
jeRFBH3d89G4EsV1ptV6oGZ8ADWtoccUK+6StZwAz3KQTNw5JcUWyCgf9hXcrxjAFMIQs0KWIoPS
j1e6df6j1Oqe9FI+pui/rycSVyvoxEN8qNqQ6QHCi1dhTz6wJKJsI5jPVyb51uKZ8/8Dh+Dme/2D
51gq6ZWNvISOR38UbMHt98A4T0ivN+i7BXSNznfxNOn3UpxTLibloHht31DuNPhduVLxXKCfbn+O
P3oGjI7aCympks3D0tRw+50m8H/RpomhznOPTYo10eL7FH1qOfQr4ib3uWwtNPDU9o0sW6kdxpd+
k91tMbhYm6EC5Peg+R8tfPq6fxi5+pGkty9sY6U6IZBK9bSG6/ewlLUdqeSUXgukyjtCSHWPqpVg
o0bsZH8HyjeYRcu51PuxlJP/v854iP32HtJ5K2seGUxnEhX0nYsf3dKfz34QcoioYfJHnWtKvail
63GrJ/uK4N3wpWwnxQFQTPToFgvO2a+aMsN7RPf4szM6Bn/lGk0jF0DF8X4LuHJDkfa0cmb/u2dM
HPqfS8bi20fkJhVK0obykrIGn0aClBFaejRVkkpDsVcx+O7xhhYOxoJtT9E+vm8MpQddn6XsDgoL
fpgBpWaclFRBdVZAdpPfNZU/9YmOHVyFOwwNfxfGR3zijGjny2Za3hVDwmmwz1+3yXVeZxuW+ETS
XIbiNxL9zX/KHc6uxNZ48So2JXU6L9bTQBNX2sGFLtKB43Z1iJ+SWy5tZO8AXWW6Uyf/9FTDCEjQ
RtZKKqmtfAxKFfuohhCJuKYXJfsS+ZxSMOHbcvxAWpR/+rJUHfZFzRTo9AwvUghI49ET8PmssUwL
D4M142MkMJeq5pZdkiLLalTUs3kTrfHDCSUmeY/hvb4l28OKqNAuhLrEv0psDyF9AQi4Nvl7fAha
WUxr0OsURJODie/HDxDT0Pfd74z3WWb6AUo2YXXK+kyJikb3u57DH53xXLfoqKXCoOFRyalnPfuV
7k7b2w9tNHXjt/g7UaIETuDBn0xso+tO4OnZxtpxM+HMJc/LPcOM3janUAiWyEdcxEO2NQcwfh6+
YP8deVcxex+cTlPE3Hl2066NYrnrFPCsWoZ4gG6oSRTxiVUygsBp5/A2sbr+jCes2p9CtKtmR/2/
16mBU3tLHX3DzfsubIQFltmErJAxgJ+gKuMcs/mzE0IBK61htop4xnHluBnUKdr6Olei0eQBFOCm
QxX29cUT+DcRAYv1Rzp9D/eO33fyaRCOnRuZw+dBnRnwER3xnCIr7Dat/AuQWa5PxpR9uLcd2Pjc
GcQiCraWiHMAz4pvTRp4AE46u94Hrwq8q96u2nMKg6F0Bq/Sq2gzLxoIrmXATU6QGpyDmDmFXH4M
cxx0iqbunAKVlsxCL+4sqfgjhoWFD8HmFdx8B/d94xjNAP9Fzuw+tANH/DMTrJA4MYyt9V7xSS89
Ao5AQg9PC7RFIocVKIy2u/IQjNQsnRffHqSP4RN5xgtc92SVQBe6iPwxaJAP8jzTRiDmoYZi0Nkz
sGWTaaV/E/A4golyaerBUXH9CuTn9gRDvfZX2evr3lLbV3duCSg3jeriK3NdESqnK07A/4bjqJt5
C//DZvByuEMMaoZ5bOku7TEVdj4oGoKIkkNo5uwhsfyMtA60sJijsd5FBf8QKVAZPRJtVJOIFq+b
XaPgkNQ5V3SSbSm1vVqdLlkJM9s5xxYIqxVv7I3wDKULXq9tB29oQXu1pt57SvZwkbUs2NjvjugQ
xALhj4/vurC8PRmod9DzV4Bsz1UmVTnVDHiPzwHAgn9uY1+nJqIMfFcEuU7tdOMg7SIyNiMyOEJX
3Jwo1cPbt3TD6GbRFUOvyW2WrnyhMrt/O3RbbZ7/vIsOPyaqAYR7w/TWWASF6BqMq1QmWI9btca7
QM61sztg1ltR456WveCDax28p/6xVgvhWlhYAqioSOj6wmFORMKTwiOnwSoJ61ClDCfKeqkp93PV
XIlXOV8n+lpatuWL5QDsY36f79tt4uMzVhMQBo19Y7SLV5ueBXASowk78Df5itftfGp7up9fR253
7Cy/l25r35cSZ2L5knockmkogCd0Vu2FHZ3MBqfTsNj0rikvtveGnoNeYcN64kdoX0TshpLe1//b
C+lRKrWjDtHfYsKFOht6TuPgKV5cWa0u4v4TTSVkiu9Mt+c1B8nr/AyDYl6bn7TxFS2P5CxNAaHI
OD2QyfVA3K3BAkMUd9x9eOisxnhnatyy9qJ2nrSPvpZAuEScMr70Nb+yrSxQ+Zk8LPplTlYb1NRR
nEvz68uyGAK/rneo/bKQ1lUgTVVSGu9k3VUOLxJDEso6Sw9VwTgmZn/wj34d6yTALD5uHp3qhZSu
uWf+ajjcfKA1Jxhsrr1R+oHpXe2I51XlkydNRi+/NJtcpYTjgR0A8grAVZfm7UcR5dj1L+/QIHl2
kscyNAbL4zdG2SqVZ6GOVtbWcqS29Y24+IsF/zr4TVlqiAOBYP2yFqMgAE/udn9R96cG6KUPmVLv
yfQwlCmNhEk4KWXsFcO+7WMl1+tPX0/1MR3Ob65hvpKNz6tHrot2laE3TU/LB4UlJyVXW5Bwk6fp
e/kuyLr7RepVpl6izMcpbtaOyte7LTEKDMjA8zu2hYx+Ej9s4lBrwjOPGS0JWI/w/chqfWqdgRrY
8RA7CWwZbSsgyBcExDkRLDH4LocUfoChRHMnGBqzYf6WrMCswhaK1oGDgGeqtiAw1scYvG3OxWZM
I+JWBZ+geGOITJZPxjNptcPujuVSCtsy/ZmQPxgfPxG4qLk+A8gqz/tGCUTdzsL1EAG5tGeUkan2
kwRNJHx6NkIMs8W/nAjSLj4lyd4niC0WI13PXQ+u9r8cwLdy9bU4SYa6x5R1ix1tkVoPNoujnW8W
BmSxjCuoh9CvLpY1bgfTMY+i24Hdhh4dpV8t5Xd/B4Pf44iBS+6UkAvQAshzL9ZsLjO0BVGvCGYz
yWNiOH1m5+Sf+LJ6ugiRyBnrN6MQPAWLVPOnOGfEMeZoihS4jIR1xdUXsWfbi+o3yKmzZ+A5F9lG
pW1sP9T2cN+5TsAEFu0Vt5zmBqlc7E/A2oJTJ9EPKSO9uMSlsYW75YGDsqv8YESlmz1COl+h/8AQ
82EPyzkTx/sGmzudbiCrKvogavKO9H5Rpss+sCjBtAOJoHya3pPkMFjF1GcsYDjgkxfkvp4mQvij
IY/2aBgSZN19dtix81ga5Oc8I+xX6o/R/wA61lZpxnYM08/nP1vSgvlTDI14YJSZkAMzphwu4KZZ
bvGJa3mPAdD8v0Q1g9h17Dsp2l1dRk8w7q0pU6bWOSY+dgXtPIneg4T2Ljdwf0UwPo1zdHY+gCWN
K4S1+FTj3H7ICei+F98d6BOLp6vfkYrEhHZr+NmGg7uKixEETuJT7RINNcK6A0FBw5wzU2gYR8DB
nXEvzlIJAEG2MnJuyCU/US76lT/LX7vmJRAK85Aam9zbM/Shqb2jS842OH+qHj0/qe3LhNRa8jsr
709mJJbimW3hdBW8oiDXSIXY+TXV3ya18/yWzAzGJnv7JiRfvEwQTnYKZoPE1W6Ig3t0qvN9HT10
Ex20GBCyHKT3ifObjsGaGza7HPm+PncxdZHgOZW8l+2S7HAsKPZqpG/rpx6eFnlYrWO9n9DYi70O
UU3V3kE97OePG8P00on+mdhBXMwMAJ8Jr1lmz0fR4I6aDAymnYZqXpVdugXm7ars5+Ylm/E/zqzw
l00DKni3yDuGkhGcpIz/7PuFRSGZan8OU3xL9KMWk1pdSDJd0q3Z5/J36YHyUAmxZxAD2HINnVyu
FjaWEtWoEm7j8TGzrwLyx09cAfiAKE6bChBDvDgQKGroal45zH4lt7F17u/pVwbRUfBgVrPxepEi
wGHvGy25a04i446H0F44y3Ph6sNIvyQQltK0yMVH1ELaL8lM2Wrq2kq4OMz2rXwbevJX3r/6VSt9
qO8r7lwo8tkhUxTUFunA/g8lxzyMPFdBcXoyS/9Tocqp1+CEb4D79QaDnmo+UCcUWxIDc8SqXD85
EkHrz4kTZCwZN40vMs19Ir8mWIITzsX/wvWFp7RurkynhSVzx1FlWcXI5LxWuJzzhRcE2vjtlaXB
w2T4a2Bh6KAJ59ziSwuKcX/yO/pTjefPMrnKcZg5GDPVBJKSxBwmjOmd5cKF+0MBmAcF5m4VzwEb
VDXd228OHP4QbEJ7tYv6Yne/jRjgOANGksKiLjhPAtmOKH2DhMBYFIOqdqe63c1RhIgrUffxAve2
bTJLhaLb9dDSsRU3/APNr4Zfp7NoVBdq0c6ndASiFHSWDxPefyvNr/ns0Uz6nXq1MsrVeKKqp942
kycCqo2O+NRPeV+PBrQ/W8lGS40EReXLjR7XWWq2AvZHCDzC3z6ph49c4sVgbMuPk0BtoN3ecnMm
7oTmAJrFr8SCKGix0h47vYRFmkkzesFtxws44JrnXuQvKuM1zM0iMTSAefGvmr1COi+kJo1pGl+z
Xl9F6pv5qe7VW9sUuOxa6fCGX41hOjPytFfyBSpBKRDNdbuzDjn2iX5kZh1C32Gug0zA91G863XT
X9VSb9/bZmOmniCoZgeeO+b/QsoE5q2J32DLSgvJt+fDPi/CVOWSjf2iy9oANlWB51VhCGR1NGQn
PnWvEnxuamCIaCjPpFPymiZFFdbiSmXp77xR6fN5VR43fDXb5LwUC03FNhH40ZtZ7wLNKWADuJv6
CHQB2kh8HVmmv6atzsBBJavc9VztrG4MA1NR8LHpEmqTS+hIfZXlwlh7z6TKnUSppym0H2ZM12Ez
6oJGs0AYECduRiwLgXgvE7WbY3b/lBLEFo/Z3vwAZVPmnueWWco8xNvFB+Pt1hLN6rEogABgFGx7
LaUMTz8EGoL49O+5G+SHGZ9xoQzNIvuhki65ePrgelc9dnq/rlvuIeN4uvv6G7p0kt666VVEN9uc
2E7Dx/BIOvYDwwsICUJ/rWTkbZFg3l/D7MvT8s1xBD8BjBJVjdV2Cve1LEoiRpVItB7IPe755dfi
A2cGSSWemG56OPwPnMgjBRpnoaMNXeZlf/ovAffxs7SOjPPkmb6l4mv6KP4DNbFey5BplpHaMsDF
VGmCm5g/z36xKglgQhFaqOhwUWUAZ2E4fvKSwKHG0pJsTfa3ykamnfW1GXmxYQ0hpqoaRq+Cjo2W
CFZYsL0jbswZyV1ewohmawSpcbsQGCyh/kCXir7nSVKgOaV51zSUsAXVCVXcj/jiiA8bFNerC6+J
dtPk/ZkmjcR9T9UCR69RaDzm0LD7NjROpX2GIp4d/D0LfpTGy0cFJhC8BPbu95At3aqjRWL3xKAQ
1aei9cuk/k/5Oe75d4R6506jmntFz2JZxxT3YcHJ5SaCg2Spkg98UA4kjI8kxpnWkYo1UZfXQ6BG
b4w6Hbbc6L0y2IeRX646YK3SpinsCO1LjM/2wSRa6Psq6k+DF0EBIoGeiJWB/36rkliEN4HokyHY
s4yJ7MHYFMgAyV3Vy0wPHLaCn+mVu6gUftD7U/8ZrVeMG46DqSbxQSVZvr5XJKEn81kZI0Ba3tuf
J8MIatiFTssNhs70EskM4JLToVCyZuIvLlLEtAfW5b9i2MjVy8JDfAwVxH+TLZkSyoINfDDwfUJq
Y3ety0bRVomaJhsqv0yFTtEAz+eRmoTVmeQX/Odc9fG4auzzwuQRRey4G7MXeTGf294ysME3ncdn
9YpbJ/h336cpzMbR3WHPcyjCxqBVnTTEg5TtRU1TDjJxUTvTLxxyRNdv/2mDKYaxR4gKJD6e1Cf4
PxMs3msaGPOgBUEBEYdtPfN8S9SbSYh/ZnXwIl3qjseqDa/mt2XiXRmAacvSTVsUCTCr8jo2OkeX
sijdimV35SMkXI3YjAh2JS6pOYQvrivXiGmFNmvSS72yPYeGUptRyJZBCGt6LD/Kmd0cPrVBcl4q
jcQ8Ws8CoTzFtSTNVIrXrgB84wt15ANOOkIGzSmTBZSsXxg5I+sTOfz/o4713ySqOusp+XaZi3ZO
WUE9oByTLcYQxFU16n0EIkhod6W3eOZG39jHUoaXi395bU5HkdTl6pqZi6nNDqIFyXl+Becxg0cR
5Obas0w08QmdIZJOfK8drP93084NdjelGneA8GcfN5MIM3RbNRqsvDw2vft/kYyhvz0T9QprBbWB
W87lrChd2FQuTLycybsbYf480yJ7kxVmxR9X1rms8u4HRZ68R9H3KaHZHYXU1Tv7SMN8rcioFFlV
rFtuVt8bvCd+KUKpWekJbc+Rvsq3Xg5xrXvhsGv+jf1JgCXXuFqILK7MHr5ZYlhQuxUE1+185+Y6
aYmc8Kh4kRDVoyVOHLpSoHIF1YAXTtwTDd4AEyMeAOu0gzcgLQq1KQj6oGabzBJkQzAsLpv9s7hm
sUop3M2jUhT+JoomvQ+7AiAxTxOxj5JSvhIhtrXFNHAXDEW+Mv6tBhx81clX1LKkh9YRE6mlj5qd
R1SHlLwKIUPL+hUyvMJAJvNdUixmJJdqvR90J+cuj/tWtBr/Fp79EioTuj0tNPx0xpEkznVZod8X
Z/ZMhJwaPYpTujD/zKievNXXsDfbUgX/SHQG3zyZc+F0pzcPCivRiPnpxwq8baC/6YNJcxe6GweC
GuPS0rEGU3Kt2M9kkxeofI2IAQUp+9uSukW2mbxsQ8cZjCfA+dHAds8eO4S6KSDILOFczKQ0Q4N0
gLIHbArLoqhvPZck4aQdbzufdNDm1bn2hGBG6NLTm4FiMjgRk/FKCD4DT5CXGRnMqOvIX9XmlOE9
dLhfnYoyArZAVtAwVGCk92wNNwVkvne0RNgjLymTMuMT4QLLPZ/8Z3pqtdHCSHQgF15I9EYghQXb
8ktqWdgdmPoXhyUJ9m4tYGXS/BhiS9eInC47Fk0T00GDNf6mkXXtwdTvNdiLX8GhPt2K49ALC9x9
r5VVRaaRV6SnEKXTo4REKPNcD5SLe12tulwdxUsZ6O9aJmou00qan/78gWhAGlNyoCLVnOfqRgan
E3UxMcvoirhj0gy4/e7myJrBhC/4ynsSomywR6b3kLEyP3PLIA8C7ZBPceMiBso27omhdHdGNOMD
/TcIThj+KirxtY+Yq4cJpbsOpOtgDYPLD7ZY2AQJE3L2Xq0kHnt6Ycvj+tnCVI6LyrCdkNytGf+a
WUoJ7eM2jZSGKaA2bvxNHFnV6lLF+47OHL0Le0VC7PjX9l9gbdGyW3EDo15Mn4SxSdpC18ZCNtOK
5LwQ3GpA2vZzt3CQeT5G99JOO5xI1/qYqNcjIZmNGb/h+gexQNfE18N//wsQQqNpFIJ8viDw3pKu
NNxpUPO5AvJuw7MzbDFP92bvdb3YgUS86UYQqO+e/EH/cl+6VsbkoTG4Aw90T1Kp7vz94zd0zq6I
/zO+dLWf3VFVErPX164JAU/LwXGGQcUqp9fgCOgdAs16vyUr4HWn+Uwhp4H2LYSxMuu9hp+bJKNI
JKO2PQknMVwcTD+8CI2o2ILBSdbKo8la7GItHxcbVxPCTt6lWZeGAm+57a7PW/59TXGGJqy2H7GG
r0RiC8BarfoEqdYoKUIR5lJXp/aor4q0/atWazzP/Dey0tazU6PVapae4cWwIoiWr7SaFpppeFHB
Lu44cwMydLtFPBSRYL2RfgDKPliCm1RaGrO0QsqaAAGD1YQLi0o7A/P2dpJYU/P6MTqT+JqeowD0
2//MgJ18xR7oxE9GkE07jBcUcKvyawTm3MA9KlyVXukncrtKnnEGB2k88AI/2GhnPQLX2Y7MjlL+
Wa7eMFMoXLQ5ghjoYb7+OO+6PRqzAaiX2hpLoxVA5AAjoQmh7dK15sGA2H/rKXOpCdoZQsZc8MQi
geBXcj/lykr21PopoWwVZttU87qr563qIMmnjtGg6CdVjRPn4B3cMbIKcwi8MrwsJS2r0D9GWlRR
Rt7pL/cjSoUDfXFikrVkUPNgnIymOnYTw9546peNWKkiq3qHdYzls5hrIXKiwzdwjBqBSjgCgXlr
65bPexqsgVyVBEw2GbdtgthdEYLDHd7jJ98InOUPL31xj8RUiSksVOQ4FKRZi1Rro0Mce8fBECJf
14M0Vjo1njkE+NSyIvS06EUPQaQ9WrLCsZ+Kry17WfQ+cpvnES86vPgH9JaU/IRaWoTuEpb8UTYR
BOtqx0wm9s73jM4cjXDmSkQ3v87v7WBLqAwGmr8kC+IeoXBFkXYTVQCtDsEuvb6nKuQbLj4W+JcF
h0/fVxtKEPMU/a2pCF5ttZLzTYJpZeNiQ4WDSzza7euCoXRe4/jXIYfGQ/EE0hOOw8H3fOWc1GBZ
LW3GKmVcArklv0lAhGuqQQwCwwysZXmo/j36N5UqokXHatlxhTL0oWHlADYEFdowZazubZr636r3
TmmGQ6g2xhP2/52eHu1VAq/jVN+HJfnXTT68hGyqF5s6gFGcRSQIlCSjESZ/oBRDNthuB/XFY9vq
1XtTCRMOUmaesRQEFJol9Q6eo/64DMrkeCBTkaJg+Y/9fAemJucIv0a6YJFLnBh1jnkZK6ogx8QS
/7ygXpXbUAOQNCWEQ2CU46pf7LSirCI97qNd41chpVNGQf7zw0s9pDP4yPQB5Y9qTFqi3UutWH7T
H8cNtqU0AXzlGKvKsjN1WReMhLBsEXsddGK9GyJAZmzJhYbYDCsj8GeZoXoaKmxf9r/dnbopNN/2
+t0SdeBO6G+leVy5ktyob2Y2WTs9MbYwrfQU+2tVcdUSdokbMUVGIDdEdEm7af0mVjrAx9LqX+Q0
DEYTQTouf/7BPQgc7Zv/eNWpJtZ9OZUpEijJcUUvwVhSbw2ON7fhBwdVZTLq+ZRg+HLbKsxt7ffp
22xPhlIlEVFU2fx/T64/28bQC6Zz8upANNO8iuFK3M1PMqBnOvPEs43V7mhRe7iH0zGFPS4f20hC
kNwTxh3kmE1GbgRrTN1IWY9uJ0bSGfEV7GEWpLGUe7YLCAqbVk4v2hi7SqQPzswsoo+LKsOmN8h0
bK62CgGoEAOIOwMjjKJ+aKk3ZE/4+hO/btPOj29xECm1qUV02jn/v/wXYlz3ouhiKoJGY+bwlHUY
IMxiMNXVQ54OIu5+aYjxsvuqmmFcxLh2EUrN2C0ffzSeEH15G+YqOVw0j6REmGzihaPKhgUCynDR
FsVOpAaf4JZQ/PbNFlVs/qIw3pD0GutbmcXPlyAZqxGdfba7h4Fr47ubl8heXw70SAxdXhLRU1dT
9/5dnZsjPMnLFvS13WQvA7KshrgpRXLtU3aXnCF7oJ5p7rZtHdbBhkoHIiRfzi6vrXFEgQ+qrujc
kMUsFWPrrL26HmsrItNaZHtKhKYahmQoTgbQFOIVnF/iNb9UPRf1FYn4rAR9EKCWpUfO3DKqfZ/R
7nlaOnMrN9tJZ4cqkTwlp24gArHq+6UI1xRVkDgoHYrjJ0B6koRiJu85uglvB3RD+ogjY5C0i3ZT
oXCmbZUWYKEzNjQQkhreGJsH7uC6WjABK1SJMAaSDi3OIZ55CiOkYkyxV6M4IYbFPbToXvRAgs0F
QuJB9Js/ZRLWLF28Un/DocA7JC0HwN20+2hpcw71itViFSnMObPAOHiuJwvjhHp3fziV1SR2hjcE
9lZc7HOXPLXnN89evfTm+JWgCH1LsJbH/gOk3Ua2jE4cUeIneMzZ0bJuTYDHnDQwJgGIglltpbGv
KlVvn1DOmp0W/QxSF9Bk+MGg9lIqfk6X8bxzTl3SIqw/OYORm1WxfyGX1THkFD94RuhxBZwDrVIf
bAtgPbpfg3Ykubl61ZYBy8xFyxR1s6PaUSN/YHZUmql2IDAOlz+w+gm+uog7G5hxItNuq2H/dcGS
87DGkgCaXOb9+pf+TiRf3CAFJF4Gjs+4H2bZaa1QbTaN0rPfy6VcvETBP5SOCbtcHcCJPT6Jn08b
q8h5YRF5YbSsk67kjdxGjvJTgVG8yXgQwIqH4gT5qxQCN+okGrAVO7cJTjjXAsjRcDgIfJAAqD3I
cp3a41AcP2RJVpspcqbr65T9d2f1izJTTA4PuWWlOPwDZecxEElq8+Lx1CsmChyOxvgUj1K1fWxJ
x13hN+Be7BHomURp/vrM60LATobasaLvaxe+ypebGU8/14R4+ZItd7EDEq60Oi/V29qmS/PjK6gy
cJhsHcMDUB8/F5tI5aCabn9LY6zEMfXS7b8cBUPEeC6Ue6xTDi49122VtSBGLJ+1sF3eAhyfbTcP
25R6/IQ0MyLKi9g24EKwaQync76vjPbxdmZN0kaiQUNKsnHprmMCcVGqWwrqPEP3zwUFL33X+3SJ
CVaDyWsp5+vsJwLLt1IlJ6smEgczAeZI5K9e4kmBQ2BVIyHA9n7DLLkFvUxyQZcGR0YTZMK9mpCA
O1h0+7J7eCVO7umkktamucS4R62mW0nlbaT6enG75bCWvYdxN3MRx6I4r2CJRHUy6D4GFudo+/y4
3n74n6TyaQKYYYAdKmNXG432u7QPc8iN9i5nAr54NbwYs+c3VGHFAeKep9UlJe2y9LrzLzJ1p/E5
ppTvqSbQ/w2jKq+0DgzvDgaN1koFibxWHpJXuZ2E8/UYqFJYQogh23sBgyk5g9HHQzJEViiANNZ3
1K90YUjEzHzM/ojWQinbdGB92MRZ3lfctvYh5SLZan/On65ey9bFMp+kD59s1cNLqNF78/omilo7
KOEJMfs+z86hsUTr5KWhM+peYHCQR69cvgrNfZD84YCPXq+3ilo3gC4AeajQy668p8IuCXYpUaF1
oEKV1qnqCPm7+mz3+CKdKWjQg2FE1qReKOGN9nK7hm30B1jbax33wZqR5ijqbjpbCyt+yyslwWf4
l8JHK5r+RgkC+2W/t8UPQa4nbamhvxJ3ifO2y8UHaYYoalZ/10tLXnpEU/JSQLnTswMToXtUKx2g
gKp4X6oferzhLMfikvacEqb4Q9qUnR9m/QItdT7C3eMgsOHdXjWzycBiGkzxQWI7TMvix4rll618
9kvwThwlQMKKOq6tClBbbag2NEoCLk0IIMgiVxezP5FqF4JD/W9m0BbAWE3UFEQRW+Q9aeNlhFUe
KXfwg6jr4n0Tvsr4AxwQUHvdvxMzh5Q560nVVPp+RkkbBlcKKrZl0ZcuKixnWydYUqVrgFGZc29I
iG8MEcXjlqdWUiKUAGpe6TxP6LQhMuXN/3vlfNJ2fTj1Y4yRwrt4SpDnznxPoaP1j0rA1VcMXn/5
NrAhZ13JRo0VdEwNYRY9evVDJfX92mblpbyrJ5uARrhwxCZm+H/lJkjoklZZVM9mokBj/pyNYA45
5fu9La7KQ4k/wCMU0jeroWiXwU+EWKi+u45s7hqSJwH2871M+vnkVEq2HMwhS3NBdY+9NIQ8QLCv
OC1FhXdggGu4QDlqz4HAitq0jm1f6f6STB0DSlzdUdvQmEfCnpVQDYP1SWCADiaqb/1L33riTRHd
JGMn6Wd/z8rt86IydTfVqhVvKE4E5S6roTdK8Yn+k04ZU83SDrL9iWA46vP5mYvN2Tvewg9iEAQM
2DRDT9UQo1Zw0XOc4Z6/YVRqNKQf70owia86SCacb9hyxFEyhDwiUbzVkSkT4A4GeXS3M8rKsQVT
SL8VOmJW0f6JCNkG7UC7FOEdSDKi5LWiyIuCaTBYsj99rnv9BPSyBtSgqb7lWNc0MNpbFDJFOk5A
j9jfCasJSJItYaDIuqIzyoga2WUb1D0Y6DB1YPTRTt0+ccZ3XyWtuyLDBnk7t5oH3HE8yLH5b00b
bSZU1FJlvXzLhgy4Gx9gMjgoO0M7xU63xlB5v/ag0IM+yZ2irlSNGWScaZG2LgPA/K+BbHnByPzM
qxKCqnjXAy0ZypHoTfLUZ1LwtHYbWGaNfN1klcxMUbG+LBhFybl0JBr6PjMb+tuv+3Y3JlzIpkao
9mJlrSjDbEukn2ez1VSGWPxZ6e2Sdu8bd97NPxA5Au76swaoDZUvd2958iAenayKZ+5MABu+eAMH
ms8cuSRjY+P/KtKN+SSvgd2Zqa25tkOTcHMs8Kch9SGd4huosbZUgwgohrjTSBa6ICJ5r8FLYpHX
X8iqcR5RjWRpzz3vHZ6BnVgwWTryw3RVyRzjO33na/Jj2KKpzCETDS8QRx2/CiEmhxALOsGmCrA2
kx+E0x9jak1cuCQw4ntSS4r1YeDi6ehD8o8Wx/fl4jpBIg+OevHUTbPKutPQoNmPwB2Vz1GqlkLs
UVc1jYQjZ8OIols/i/315meEkeXOxYCFMTlhPZ6cfiVnDl57oYwz0yS2LaD6E+oMftu6AKMDC/Lz
pI6AWy7stM2bmJ3SCbbvF10iMlGbfj9d+If20doVXZ8/77IpLkL4Snw0+PAXgIlFxexTMZke9N7p
821Budv6IADH1ebi35TKCWzpetlK4pGSrA15TGDV2CfI3ApimN1YYHsETaubNTMvyEFNBwhOGjLm
NJtoSzepuO0hL59FWdfRXpRUcdfDCPl1j2GrMbOND9AW/ZzBeKt/a48Fmtgaf11CV1loGW73Hjgm
9In4xLR9GCDoInRrWiNpNjN/NyMSSIaUyUCloCrYcAWAYRkqfQjCrI0kYDlU8LAu4XIDbJq4x64D
E66yHFAZXqknv1aK6dqm3XEDRNADtlXNxT9UXiqZSIW5Atr7LczF/0daTgTw+C22i/K8WZXfD+lO
vzaccCrSGDSceco1N7HOvxGGJZjvfpaZpbA4oNF4BNtXEcoR9jJ5nEEOyyZYcr3QKi292d/06uHE
DgXENtBq5vNFk82xZ159etCk3d4p8jXuPuhPwbPfkRF3NddBjznPh402s4M6FipBCrifvThi1eS8
Ct8ao3I34185gMuTPA/YgySKz3Qoprlgbqp6KDaNoD8Wv+eIdnpLW5IAr9LD0pwWhgbf7LHSp62C
xSjE1FkxK/wL5W6udzgUi1GrnZJIT2+8EORew9DpFeAt095bmlZmqVjCHLxVNfelL6LU9rJRkjwf
Q138UUQ283fnG8YPF9H7lQhwxiPVSmGvM48aw8eKu+46kCjxxTximSgsMW7+/9pWRBWJZyNhzuoM
o6dM+UvzKkW1yN8VrDt3PESDDJXqxmIJSRj4yiWpMzQYLwgARNfqv4zYEPddEJMPa67HN0sN8A+Z
aA0O5WrKBjndrwbk2y1fhaCBqD7Ke4n75hCU5lBeSD7XSgcLAUrbZXw2E+lurJf869uCnPSnqOLb
MPSBiJ2IYlr5NhmUtKp5Aiyr3R0wLNP0JXdjS1gun20Z9jyswxsS63pCS420zoB5qiG8q+eUT+80
OxS/XQGr8xAFCoRQbwA3DR2qJmjkZGdO21KGKph4j8PlsZd5JDuTE21NmFFipluVFSoZI6LZrnXz
mJPhINAOuz+9K2Lj/sdJzISEW9EWn4w2RPJvJONKdfyeEnHvNp32z+qi7OMFZenHgbdEXiePv27j
S4AyCN+PkUmiaaU0JyI8NUojUnjHVEnEZB1AVEYi+g5VrSYt+P5eusTvXzCbabRVjxNVm5F5qu1p
3ScFvgGwVlo8oF2bxG6a5f/nJzkEM88trFXZRUhGHvpvDDkshwf8Stek0TMhZjsHBXqw2W35tnwh
sDzUcxyOk2Ge8wfv2Exw5/JPL4PM/49nKcUlOWTtJTo8KIRRhpUZtiezf/aYhoA4ap66vsTqkIsp
nVnuHWXiCdhDYikC1ctY8WCUCcz1cHi1z/9CF4birfl30ZpZYKeAQ/l8AwC6EAX5mMAGhheiwnF+
NyNUHJbILPYOtMtonyhBgTziF3gf5IJueDQnII3VOKO7EAEb/QXWi4E36DKqknheqxR6u94t5epK
+MNqMH5KkV0+7t85BIwiJ4l5cDqJi0wO/P24jNOkAZjHwzmCScV+TK9R1D3MzK9Ioq2Lli9Wn/Ah
EdoAaEpqo3lW8hWGm4SHFg9ImB3S2e8dVL+ebRbjJ5f3kwdh/tZkSirDan29vpBZrPxA5c3l33UT
xHLeIb4blBL1FGZPW22KIn/6N28rAL8+emi5XU+LudQsJbIxYCerL6Rf49uqRQpheTrHx1peBimL
GvV4QH6FYpO3tpQBOF6qKUYqM6UtxtBysZ65lGBPc7YRvk0d/fs16uUeyONnHtVz5NyHAcllCu4L
kT1kafsI77Yqzo9NKleAL0lR17xQpo+KUzDL9a5VeIn/J7/XM8IS9RjlzZOwQfLUSCnqhhIyxr5y
Eb/O8jiawf5hjplQm71ptJT0+Ajf1QSR0ID9RnxvOyYs40Kf+3a63hS5wy2I/wrX6UqdXjOUddiH
u1hPhpwM+He/fzjq7NTnwysCOcSE41A49zne1bL7OxmRD+gckzj+XRPxNrMFrcJKSaBAit5cmHVu
pNBmtMsy+e6oTHZUVkFLKQn1vo/T3bDTTxJYi7ACF/QaA9Icz0LfLzSlirsCQUDIJxlgpM7toi6C
JnCK+UIWivZ0ujajl08VPs1NcAeBXvFH3hcrsKCR3fjPXYuf6FAZgyPxvJ6RsGLIbpJ3gplrCChn
OBX8/SIa3Xpwtk9S0fIUJgUYin8uR7sEuG/APKPKwz56vBQ8jBx/xnfl4P1O+nqzxHa9pE2xoQj6
wFO1rkqTOVaM3TIocPdEE5MRtarbYeSyVxHOr8YekdQNglN4jqs079oYhCFm0F8sSl8yxbgvnEz+
dlHJvvi/exN7Fe2SfVAO+BPKHta+gDKKr1McxLMu3ua4LyGqWOZf83nO334qIHpWkXMUEyVIgHpT
JGszMEDJEt2k9XjXvCWeHyfM8mnlyTEYvyiQtBDpuZkY/VGL4zhq8TWfnmmWsT/ShNpA56Qkr74s
wo72lhVRKC7lZ9zaRKs1xtiHsOPq2zwcljTdJ2fDpXUAX5XGjhw4Zom3d723/EozE7546cT22vOg
D4eEeLQMdBZNrZ7J9Z/UcoZe9o83uu6kWzKCvWeyYrOsb0N6z5o55hlDaKa06Jp+2g54uefiDBbG
fcE4Yc3/uE5frexnmgFgQcXxYnuo51hQGQtNfZFATCTxmqm2d5lmE4LWVzi0X6Aj+XlJw2hK3vyG
Sfnf4kx7KuniNI46fRmOS2lE3zG4HZX93ZcW+zqIcMGI4zEfSiVtPhp6DUdS2NzRVuVcyYGqfTFJ
TJVWcc+neEFZm5CIMpBGCgEIy9d4pIdjPr4muyLNOgwjiThiWojf/SGqHjHMArWQZ4GOq8Tbhgmx
NSatsBuNbGgva+JKN+Oj9fZrPCN1rW/IDPcrvh007MABeibFlZPaeIhibCexEEH9IrqVyu5FjbI4
JA46dwf5QAZ4PcWHSLN73RQz0LPWSJVWgDADiU3+PAAZf+3Rb0a2oZLX0QomZBxOsZMomc1gHEbz
9NZd5gHYwexlgVA3M5iYBTu+d1IDHE6CUILfFnHcNiSkILsmP+dcaPQKZXhz6Glk6HhR/PTaUlXN
dHygQMHaC7G8f6mpsiwVMR88+se3ZxH5gA2EBoTM/MPqev1BoKlBRwFSHISNTa8fIFFt1tVSFa5w
Vpv8pmAawJMnWsXxkjOguAuOUIyOIoO1hqFDz6KPhBjl6lLOTBwRmPYNf/4Gob+GqtHxsrDaf6pS
T3w90uCVPYOBOdUN1d8Kaetn6zlK/Zs2axQlZIwH9L0XM5XHYqqLikJRTf13L7/DUepFEyeAWy4f
SfDoTx6dsrFHvevaNw+vq310qjUIr1P0woD3ZY4St9YNhwR8BHjkfo3CBPRgs6dk1ZTmtwhTkV7J
unNXz/05bOBcg5/dgjW1rvzuHBENNIzo9Q0VXRyWH6wQNhCTTA/M7PuvrcDKr0p7y77r+IsWT5Rf
rhUB/ZMSPGsxSU2CaOmCzxqGMYNjztilRkmkL4OBCg737/nR/CHHGMoDIjL/RTOlcQAcCvOcmZWb
UEFcP/qAeQlNfJziCCmEyn4iIIeQpNb2GP4y6ui/XmP9xfVkW51H1PyxPzaastrb8bWMa5qqQKpQ
L/l9c5SWnVqagY2cBTVJc+j4iuUNP1z7sfbZCNVWBNa1mbChl3F67sTUF/RX/7L2ST+aOlARqyur
bPAZ1oh6uZp2l2vDRpInQOnJKvUiIA8RlYxMBE5p1zfWiyryjvK2pwGLn1RR6Sr9KQtPFpNyGnli
Zdid87QShYutj5LcSZ0xU8DfThVj7jsMQQ+dKhp7qh/4VzAQzMkUlN2t6lpw2Sz1wcyzhsw2riz9
go6xICEW8/dFB14AlioVkNdnGTDLEFz+LIDmKVEbwCC1S9IscwBgej+6CJvpg2C6VOdNn8MGx5CP
EgemGyLxvIOXzKLCQ3IxgCAKHm/1aHIeCqeGwIeW1ZHRe9aLcs1JVomFkCAT/UroQFS96uLF36q4
lpeHY7cBoupxYdkMBTFgFe61DEKX4IxkUWTMkHw+XRRgF8sS9JYIKchfuxUUFfkjP/qY9tmTTQ0k
WsZHHeZJvb/sXqgicCLVdFWLtE32bQGEdNXuWVY1QHx0vDt8JVKRW4s2kXamgOBvl+WtMmzotabY
3od9V2l229A061KVy9fK9WxWHlTR+VdgBXL0cjM6BATj5h/uWiXhS3onW9uSCkLIXW/L20TsBgB9
VZmyJZcIXaTaE0QSSu1cCE5hUN5SDS4Y8RKx9avSlBQhWEyETr77IRDjzhvo/+E3uPjRFx3ZKyWE
zvYtjL66iHcgHhvjlsgPlM0SQ42OKz/6jwdJTZQ3Yoybl/P8gKz+a9GfAmw65SJwR9Dmctl94Lpy
OgSla63D6GmyIaCUoxqbmJHLYLEkjlr3j1diJEyfVWNirZAlGjuV0Q/lwSalNl8rx+qKwdZHVu7p
X/bV96KiGRk6z9xsvCPBUlw4uniy9fXgIV5nA645d5fWvJvYwU9Uc5qrigHjfAlOWlkIckqYjf/O
pPQCRJriIr+XRv1Z3IVJPyHEFb9SjUm8n2HSzJIaN1OMq/zrA1Jv12Kt06CkkzJp/20XKUkPstxd
1BSU4JxivIkQbQS/daO5E/pYV34JddLZJSfvf+TOQNmZ6cIkvL4njJ9nCr4tv6f2DofmOAlC7xHR
/K1nKf6KLqXv+fxh4aP67TPEdgbVJ1nuyrYdf6BCi+x5UdSrmwoc55kuvauq5l0elSGmUNlT2cgx
bMRIHgzaV0jzfjyb3h5f1Q2DQsy5Lp7NDjqZRq34STOki7y4N2qRbObK3Nn/b43hJJz/7zbTBXpG
uWk+A/zSRQz4M4+19q8qALs5PppyL/w5XjBW6hAhmK+IrMPJEmXDswc0hkQsk6kGM5QzbZDZI+aM
xz3cnUF/QYFQINOFgzIqkE2m3rkAI9m67q4FSQDj1mv3KBMnlvChyxHwMW5vBzmI9nvPiccX5niN
oenifQQ6fq3qcC3eT69HVUfpNHnDEROev+zqwpvBTMVLFIhn1tlIYeXgX73z8xWv7iXhpUSgawKm
JuMMfET8RF7kIoht9HtCsPSj4vutxQX9I8CzsgzoFKEMiD4+zjaois0HTh6a4UXrwLZTW32Q5t0o
PjHzHIrSS44TeI5Fww9gr4nZGhwmUfSzBr8TkS+VsKB4Vu57gEx/sycE/683hSCPocDjw/oMUoOL
D/0OlR6ACUffyqVBBJ+lb7t2GVQJ9qMJFXj0CJ3c4Um1DI5AB2WtBDkh/EYPp2csge4P7wkNRUw2
GRovlAWocdytR6TspO92oTVOKWa9ABZEIHSGjQ388We2Q+5Z35u8Gf/1cgToS2RAX5Ydxh+q/TCF
nkrMjfP9M8Tqt0tCIcMWN7pZmKthC4nbgApk+CF9755Xg3FWNIluFrJd5kH3je0Cc79TU5HiRO+F
DtZO2zGtZauTd2F5yDt1O6jP2FBC++QhRR4MMHDocGHH/5Cbnr/z1fao4TrNc/2XK2RzkfZ94jcu
tMWVIqSZf60W94YS9m3CuIkb3XuZXHMxBZj0/0Vw5uro7oxrogXckBXbQY73UXthpHd1/RLSQppB
dDlwmLHzLOqBb7ObD2P6aXbJtEb1uTJUphrG+hnWR2O7QTGgss0I1hCQ61SVxifkynfoIY54P4CA
RQXuKCdIefsKhv26wvkyQ/KuGgbG2sX72pYABGg76P2mxQdkswZm9zjEmuBiCPkHqV4g+LbBb9NX
bYtCpvLCijk3/zkfFY0kAmXrNWVuzKFNGgHCX7FQlb4Cy0Qi39CPykHrQ2RVC8plttf5g5/NUobX
4b3HnvRqdyqWizPvbgZcrj0+2V7/GeaeEaVQhUqSyXfgkOBi12hZ1YyKs02lBooE7GdNzLoh5Ha0
cWQaiE57e/Yl42zLZcwr50Zlhc8G6rAWrfUBMqfNOCH9FTTv83QnUh8H5oa2R5uLIUKw2iq+h/u9
j5Uv3cP+DS6OMbd8/AAHYUcrBXxBF1zkiKksQP2aXDmk+Qu3fRVum5nBxjmhWfILpBT3r/kowncb
+SztX0mUgKMJD5qh+InR4p0eFY0YPe5TTOfC7yAo7jpvBUE08v4m3d/YA4gTnr3QMauUaAvKpkH/
G0Rlol5DpCGT/gM24kqZoWz598LtQOm+ocs/C8o+plmgl1g47gn+hBDR7tW4MzY4EBcYAryniyUA
VaATzM1CFKU91TGG4wI/eV4EHZyVEAlOkKKtiBn+jibXic3vlWLiwBlcNz/55EpKHDZdQgdTXJo0
9zVqO4eWB3nDgnzf+Pc+qnnp0Yu9l8GDd/6K6ri+Efxso3iB0k+GkjK2CfRaPLQq84XUbcekRw9e
yqlKhM/MgYU3qOk5wB5WvJeo+Wh05A2LM4ZeNualShDGN7qpY1ZGqlCxOnNrMIQQC5CtSEvCdDbA
9vrh+QgQTPTnvP35aq7GPmrOeWnuD1wHqG1w4Gvua/x+QREeGbvrqO+dbfGTnTpwq2x5qkllVPel
2DlgB5anrKvw6QRGh/xUTD1w0ZPml33cG88MWuzf1Kjunlq+UIDW0XU2RGTyqW7Q7GxYGEDK9ay2
UVSTc8m1Tafe9Dm93+WDuCwAwz4BhUsBeFWdg+a45faEjdjzpRxiZHjaS1Lm2IF6ej0lDq/4Lsxa
ZDVug1/zk5IBmCiW0ysPEVDqC0pe2uUg1yRJbUk0t2ghs+PukX6HH0sYpQnNkhPeZy+yN/mTHKTO
AnloE17XJS3Lss95aj5Sex7I3gJfK3gvSOpYmaN4xzfJkThvg8iygOBRERUzPqUiZGBlAIHh/GIH
cFyapnPcQJUDncLhVJIVQ73cbKd/25BRv2voxeDDp/o0cODZWYAA9x/oPwnZo74faJcyzaDmIKwK
ig47MDBwK/BStPG4cQrkKOuEBckAB5cKiTADnAGWEABVNC/e8rX4GF6UeHrJeicaOR4KC7GCYUBA
RpUCR/+ksB75rCCH9VoO/TvXWTRIdN2vsmQTZbROqmsuh5I979hthmynUTJYQXi+Ey40+IwMGREv
qRQtDxTAZIQ9/xTxDpaXs5SjAJqoEuH2oQPMRo3vFNfr1mtZtlzQ4mjh5A97N893Sl4F2NonrwSK
W//CDUUT3XIAqIP1aC1WXyzSndbn4mwMENBvLybFAFCHbk8NjiQr6Ckn9N0cKRlu5uQXWKnlVA28
LCS9TeiJlfjFSoMt9YOEcODAOs5V0VjQZGyBpOp6U8zBgbdZd/hn5iYNjIb7w/e8BHvyJqw+F0Eu
38/0me8LV0fXTKFGMc/KDpXRsAVWJpgdBJOxvs+YN2lPpzd9E3y5iDj9uiiJrw7x/qvAtocuGLfD
EiSNzN4Ru/SOT6FPXF9xwXdelqgW7CAUKUcibfw6NszoVbegZdGwvk9qxwaH8AAMufB7N1ccLk3k
NZ+tO4mi9ac9Ns2fAHL15XEmnq+XRbr35FSP0Ab4Nb2DhO9cYGf5GXR4Nd5EmPVQB9QqjTPDj7au
87m6f6VXjX0I8eCy0bU8X2wd0pIWQhqgmtxqzAH2Ro3EH23i5No2PlkKS9zVe4bs8mX8b46o3ulz
uxx96dDYzB4D+gHFjuwjJS+Mm7LNGDHHsG9WgIMmT5P25CgRfsPO6LsjaRd8LtbzI5GatFtzZ4jP
X3W2BEpkUzJRNua1HlOsRnd3Dsk4NwEYOo3P2g6fhg6uznpA83/g45aTsT1mXbzKN/xD6LL9KRQ1
Lm2C5/ZzjZzDD9vLY3YdD/C1jJmvDuSG1T5Z1CJ+7yolkfBoWMN85br/2bfkS109KjQ5rTlInJfa
atEcz03RHEfReIDKSmwTadpmFERZxdHuGrvOHR87KpVfhQCjm8eFDWXL9NC8nKfQOxciCO6gFUry
CM9o4POm8apHfoKJbkvRaZwNshbcn3+eBGENq66wA2kCFX19dR4l5A96iCW/xKf6Ghh/Ex+M04Ra
83/SewfyJ9O+O2WhGDHFNq8F/ZwY+AVgVM6lak53TmLzfaQ1GDTe0hEf/kcelo4zjkk9LDw117s2
/3TXriupyLFzXHN+qodNeO6QfzuNI/I7Q49WVAlEjvBW/WfiDT0jgmePK6z0qSkqgazX5SOJf33s
m1Cig4evybwI2v0BBaLCkt8Hd8LMDMMsLSmctCwf4t2+fCkRVJDbspu1N+72nn6fR6fMWVD13+Q2
RiXGzNNP+aXvjtOSpc/Dvl2gdXYKNSl4Bgx+GYhLmS/RsSQGaLEwa6zJXMSH56dUgBeUGzhVzv5x
UGi/oyy1KdJrynxHHZL4ZaNjyWxnJoY4RQ+wXQBzbfsb+NFOZZTp4JDrWN56We9Jh6fW1yST2mAL
mFwsGNtYrfsU1em5afiASUGhy0BRyp5WDBQJ6Ox39YUOBuElEYhuzDEVhoewoH6EYVqCFrZZsEOn
FrWFTyzAJFIvkq7FUku+8lkLGwJATLi5frAm45Ag78we72ER0I88p5JfI0yaoGf/noqVH3MVcCl0
1xB3j++sAQs4dRQjAL3uNhLyHXQmgYwNphxpIewHgYrA006k3GT7sEw02v2/GrZIRAVazEFQOwmO
5wTiviQDTAxXoLoJOWWrpUYhzXyJx2WoLwP5IUcP+V56C//yvUFxK+lWDKu/glGAE7RGSIIIWXSq
TwFMvV6V0M0b1LHH/S5ghoiWlqOSauX2BzWNn3kdyEiMkA3TVm/KPbJGSOOk1PWfhDO8zuhV11n4
msR0vih8++WUvcdxRS9AZx1/+vTbFQ08NHN5qs2ux8JoOG4fz5chWPwMk8u8ZG8X1ShB+IlKEQjS
fELSocww6CQbZzw4K4zjw9h0IFxw/8t6qx1OKbgJ1KdLL1uQ+sUnL6BMbUk7kUouD1O7pVDOGmD1
cf2DEy+gZs7QmF3eZH2+OeqZkk02LsBY0MtKM4v3H4jQkXIRk1f7mkbjD9rpnhXHl1k5G0k+b9c8
nPVJY6v5lbovFWZ+d61MB7IRhZRrlU2zEY4maVXzwcYP17vEfiXR0fCbNkx9srjp9KcIQkoSDvZ9
Iub/hi5yZfVhHrxyZIzhSX7fyM2hgvNQQKW9Z4Nk+UfeyN/Id0uiSXS5FJ0GQ58pFXZOGZwWC5SI
pKqDfhB3koRHEQ9NouMzEkfEqckkpDQ+HYu9kRbYRLeXV1Go+qdJQJdcYgNThjAyv8C7mN8nb2/Y
vz/mejPiG38Phsy+STZA51y1wby0FhhlJ0UQe+7jfyMYibsPMEbAcYB6jI7zOPXlrEZIZ4ZeRlp3
V1GUO/AoOGYvGxlBTLBTsdi4wGQqXvQWVr9sh6nfyjgZUYFz3qUP8wRq6t0b3R3nD1BBqqZmgk55
ErgkiLOeW927vXNTyyiiQ3jdqlJhK6TJ+PUSHYULE8PSR9Rx1XlU/xeMCfzDqI8oT396SzvdO/Fi
ioJBXlijJ1XZHCqc2KvBCPM03MKmNMpxPwTsi7h9BKuZDoIsnq1VDD5lL/tgXKLN/jiZp7pDDwqX
ClzGtV1b/k0OsDtKdN/uAcxOKjHgfs+omsfPsw/IKv4IhfSUSgHP4Y+OlfflC0d+IWpPsQ20EGRR
dZrMgqcLPr+9ISOaSZopvDx95McF3tfpPgLwsYGADOV+mKDQ9Gf0KyKE0fvPTFZlfM3PvnUABkQk
sY1f2nWShtNKBEpS8FgCEWh60jU3cq9XjWN3twEZ6Twl3xxUYtlGE0zbGWglmLp27D/A2fcTyWMk
QAD5fEQCyBX/p2W/zb6kdy2VjiX1OtTBMMuWgtP7JMaLpbjjO2EXtrHX/gvebK/jxcDrUej7ca5z
uo1Ke5Kdc8xCZf4pATbOCJfG+nHxeJ6qTwrrjz8OsbkCbCOOaA80TN3PUDNrmZ/S+uyoyPXdAQ/Q
3vPtSE+Db45dgeFcT7VmnP4AsDn+ohmOnRFyXz8eIzfjHIeniXiA/Jk1DHujzKr0skOiVQm28Obu
evfNsaYdJbDqxZLkLBZnVgJ7IfVPY1ZpGJXKKoW8oQN++NEmp69s9C9pjCocVmgNhhreBfhIdVuO
3PI4WNPnBv0xjUk9DD03MAWqOuPzXC6z07i5O7SOvQ67XbmW8sstQRw9FlhA1dpmS9Yx2GsrImy6
2oAZXXcTz3BlXqeFPfrDoMO+U0jOJzbhVPMbp4teRzL9oRyxhwdWXnlKWFgs6YaajtjagFwavaO4
KVXFKDap04opMszkgzvclk3ebfz8u2+Qf9PjShdMqFkNI2JeIRT5YmAPNszWSqT2BKhA8+6vIpGx
sTNl583WtEe3NNcEmCwtEm1boZ0AzsXRLvikdhyizKMzNbwBCBW3jEU2c+ERg2WKh2G4ochPOXMD
9Zte9tAvbknOoS91fgjCynnXiC3iZcsMJXt3FaFpYarsLmqdWKRKPmge/PQ62F0w91V1+WFLUWZk
P/jJ+uv4UUQq3iyC8Te+eSP/mKBTsTcdOy45KH7mikOU5MDnEgkArAnlodYKi3UGZqRG1RO1LBia
QJO9UiYORFj3inlidLYmMvzA8F7ndaZwkT+UUW/yP/Ff2z6fdMJ7iq89RO5DEi3jAMO7PpCSwGFY
530TOruysGrflncbO/RWXFrl8g3x8iGzhd+aqUJzV1W8CVfn0nab2XLUZn7kXPpTFeHyewkHYGoG
BOXlSOYG6lYP2BAca9DPvjYfx7juIJ/JkV1RlACAmqU1rRLJISvBrtKggFRN5A7cOrOuuFC8BUYV
H0jHvTggNnDv6mVWCv7EWn7+JB6ew2BzxSTzIY+KZhebsXoPlx2q21pl4jy0x5+mdu1D0+vwB0Bt
7uMw5opGY/vHw1MJ4e4+FwTyGRZxdv32CwlBNfH13Q0nxXr7hlaJAgtgBs6hQsGF1DH5BCp9lbL7
ID+pstJPfOtfiDp4vmrRbWuzK3mOy4shEQv/+wj7smEJzGxJC4cJhk8S6TWg4WPsgNgq6TtKuFeq
W7EU+Mb3OWS34ynC9uw4KI+IenzhYNIP2FJgvUGkEWuePKx1Ea/Igyu/EXS7tK+fDUyGg8LFcPb6
gzt31DClYxz79oZXgByA9pS4yj0SQDkFf+MNBG12I7WoiwgA83xqXLii/7KZ1IGezF4L/yQnP07/
JAO5kpyiWhYfFGQ6rpSQPmmGddXSjOLFrOOS3DhyHz0cvvYSNZSbKdfkILykQDnECd0WRMvBwRVJ
5ctZeZyT6/D7uy+4OiA11fN7xGyFN/qRpaUw+aimAHsN3mz/eqks1H1qXoR4iqagFFuQXtgz302C
bKUkBL2noalctr4EKeHKP0sGyELt+DmnSHIfglihRMGcqmau2BBbZnGe1fQzcbUpghwfvTq0WBxW
XRopy43tZT+24SGr0bNOYy8eO4+9HQGt1RYVzwVURwW6iY1wNE8vceY9VukL7SkLiFXSamhjFe5j
cgSOti4mBNvro5ULm2wmnkoLSQmGkUN6KRk+s8sBFwHz3OoV+JZRR9Pl6zs9gSfCX4JrKcHEtVwD
EQG+wtnRJF7O20Z+mtworRn3/1CfFwk6rt/p/A91zVcMNgzuWsdRN2eWnmGgvJ1CFSJflhENBLCf
nsFLwTekSNdDbgswkpDSqRQNnz3ZfpEWNStv3Kg7tOXIGosDbRemJefnbJFPdyEnXddYc/nl72SX
kkcBGwIWEryPm26WlvCxMqsNKr6ozdTIJqt4w6hKWBxOCSg9OVS6fyglQPE5HRF339Qio7PAEybq
0DdPWBaCE6YKBd7A5CAlyBLAzt03sL5SDSWxyoGJnXgIjobKRBg1BLA2riz54QKiQ4vXbMtF3Gk0
eCk/HqltOhUMEGO8tk1SXLaAnQWy7CM18YsHkowmY+KODc0FDo3IWq3b9n/AXr9lW4kPloFxndLC
Ll7hBi0BJvnjvVT4pXiOfB2238FfiK1cAcX76ZlTKT3Rd7xpkZfwDV2nC+Az5r2ZlCY3oypNxZ+i
pEZw3r1nYDj3a0MnzCGKXkZgZzjsyQQIj8Jx7Fcp45AVj0dC66cVP69gopG/xANSiX9Bq65cv8K2
EQVW07NOHYQcqqFLlEaeZ9AU8eoPrKYSFr/Mga4Elj3DxBKDiMhdjCnWTxkDD2A6UkbUEYO0Fxs5
ks98o+dzeiFlP9deplz673ZD6UWcNunCjpponMLOWYgsFbr4BRhYPVXQ+VtInRvLPtRen5u1RWEw
8Ov50oRs6b0Taxd6vEvD/qQ47MZ4rjFNw4mE0Alr55YAyMoGIgZ1/g4A1sRtNYa795yIJK+KAEOQ
jOeX1zxIDWxhz6VG1yXuzycA3/cuB47A8Yh2Og4+GmlYr5MZQk3akerb1J69PLEmlI13r8UMuCS/
SrJ0cfJ82XI2d1HSxgmUID3pXBlkZmvJSQJ3L/ERMLBvLpJiwPut0z0ht9ws2G9MhPHfJDv7IWhG
NOgD05OtsK7Qa1AnwLMT0t3ir4QsnN2n7+7Jw3t3KNBLQum5pCfLmOY3FL/XfELkxxlXE8r9aAQS
Y4EqI2wPW17ta2q14Ffdxkf2pKTJA+xb4+L0o5kdfCX3UkdDSbX81FHoxm7gOkkKmJOXmCRCHrzr
xy8Z1LBg+P04Pm9LHwqw2ll/lonp10iPN1ctS9bQdfeoh4AfOhK2Ah7Y767lXGYgmksiOonzPoQS
mzajrHRm+PYDNp0t3Q+hUgNb0EtsvA1o4RBT/wq/TWZhXMLaU8NHhUcFVqy60M6qtrnZvDG63BvD
ge7qODoKLpFHytu435/uyEb0neqIOlza94zHrni8AnrGLKWAcRAsHWkWcCDTsiqe1x6rapjfpeS/
Q5kenHzwGqTYrqXzwCeYDZYzgzQG4u9CWOntH+mNJg357Xhz1uWzT00Yjmx2TqqcfdGrQFuilqyo
87EGUZ0B5RnQNwQ9uakTiwe0aRZnPCwIFZNr8UwTM2OLdtvha15bNSihiYdx/ny2kjnHqLRLPHar
qmLzW5arjuat95EcaHds8ap+NGYEuIcbT+oRraM0kc31g3btokXQlHUVkyx2OOCdZ8GFhpsuEL0u
4mto/ohy7HOEb4sFUBPEsROPpwG4w+xCJ969zd+8E7kD+SJ1UJStlRPbk7VA45wBsbG0emwpwVAV
BEDVA5MK4IkTk3MpDaoiD9fom4cGW0AGgqyM6xJK2AeLW0S+G5JTD9oV9z38+4LWDNdlGhR4KyxO
OQTxdOwMNJTCxO8JDU+O7PVBEtMQZGxCPlLKh61PyCgDteBeVKMQxSIydUveO2Bu6T7H566YNd15
NbEcwoyrsbigisjr7yjpc+E6zWrBsBVOrmDJkWl8WZsDEIwefrmuxdj+OvscwktvAwOCnRIdZzRO
6j4kdrtHdMkJ/WArWRZXN8HIiM9MLf3Cut2BLBpBzs3u3qelwIIbDpaKwg06En6PFYQtZhseDsd/
nHJPrezYoEuwy+Y/CSAfLvWj+WY72iN5u102qp+TjGFi3utLspMyVtUqnIYAPa/TaR7Iz4cLih9z
tRhFPypQbJVreG0MOjo//8zjrOUliFeRrFWpJwJxJr0EbDK+bZOUNsyl3lwHhBWM+YGPitSJ+0MZ
o8QniDR4YJHdkphkHoLCMP67ZVg16HZJutW+yR9164G/6upIfpcz2JebOgoNyNpyM2AvmwIOtcy5
8UsApcrdkQRQVhJ12Mx9oYFMfF9KmtVGQ1QLwxdvq4+BfK9Bq/0weWGRAth/7dTdiUqOlXXYO48D
6JAa0/9Z6PvT0wfhjwPQOs/KUpNaS1mi6nlKiKz7iJfM6F2wi+nPBiXTI7FGTHqFm/ARlzeay7x/
s4ActK2Lbfn0gU6K8L2wIax1JTgqNcS8Wn/l584JNJY/M4vrsoVflWIKidr8mDapHSmD5vpf7v/8
mDozSE+deJEPQvabxBSgCwbYQNMChcWS5sV/IFRSy0f6mRz1yxPqeV+4Pz0Ez6K+N7BxusUa+m43
P4/fheOiIevWBFti1MWhYRS/7UFdJlG0IQ4lyhPdWwkEWYlc1QBU3h2d0tTb6DQ82UwuqQteSSVF
Mvo9N3yykUHKTfu1XQjDCVNLItmE1qdo1dGf4/fb5OKm+4UOJDiDA/6TWnlNCBu7xrwEJFkPcUgi
o6e3w9JOYKURM/+aiyff3P3Ik0aREkdeu2bc2evm4pvn9Plyag45mYL+Nhfaq18vmQqzFPuRLGZq
PofSfDcmLHyb+UuoAWIxHNTze2cVqew5AaluRfBeOXqnHnMeWGRAGmQjyCdUOGFENiI8tg0Z7NYn
yq8rXUhh6wkRvoeGmHCed7FPctHU8aQudi/7rgHt5zGhpX35BQNoNbelHrStGngw1ifWTl6oD3Po
0YoRJFBCPN9WUpSpfvpqDcNiYEQ2LzkT/YNLFrCjRl0wmgDJpoflzCtf3Y0Cde+m8QXAsuel3DbD
zoQkNg61fc/GenS3DuNwFUqFB89dTVaNnB12Lx81LC9RcVou5Qv1HBaU/qXaffOkKFPkbMBqgpX5
eeDA9jpGfBF1NbtubWtmmzLMWwX2MI+ZpMgGc850zaXuykgh5UUGcx9AdTZkU/ihF139UTKYOPk4
6v+V35hlLMU9OBXalyw5Gmwj7JIHK/miDKrK0dvFFAuC4d8XCRB6UEsiEbgph4zEbvHiebQX0GBR
c9oYwbgXKnbPU1WClWo+KgYEc6KL/JewwTocYkEY5DWcBswdvsWvRevFhs2kgD6B8tD54FRK2eUQ
wWN+cY+4gu/VFOeEbW0jcgIuiILmVridJZcoLRxTIDUwIMnXcqu+kiYgK0X38G7wCk8OjRL6RRv3
IdnrP4aO9N7NwqKJA5clEFn6OPV7hvkZXuy6y/UtXJhp5ePAJNHDM9mOG2MvMdVcHUudKkTF6Jav
j/ZaR0QXclHiESRPYXNK6uD2KQzG0/ScuhYKl7b9uH4qscWbA9su9D1JFFym7WyFrOCcAmksRjzX
9qYBW5p+mSHq/xHU4mIMfiXXF8lqaKbFSFnnrcFiOwZj3QHYCQ5I7ZRSd9bz/HbFvhUF8RjSf3sq
J9xdjsHeo60LWXXZQbkCazSyBZiLBxMJ/tMS1tgUe4f8nzx+dzvpMVQwWwuzw2lmk1+ADa5A5MCx
xH3f11e/z1ftdo/bX6hP/op8a3sYjRUBY6sqLQlQwNtV53ZLudwvuG0sEg3HlVYkrN80iBk9wZT0
fz/vwu1NQG690uPQKDrDC0m0yf0esOFHvut+4iBzgPwLkcIfgFNVy0bds7csDBfI1oigMcW+GoDu
4tG5Sc3+epCheitCkfDJRJnkKxUTxS9ssKXIdJbzQ/d+PZppg5TJrBeD+rfoJtjllMTCTGPNt9mm
wPUXkc6G8pdtX4P57uglT/JXCzIo7slq7YcAVflDqJfb4Z7YnGMf1lJJ8S16iTDW4y1D601ko5eN
tRjgrP2HFgztsleLrIewQK4GOFwKzqGRApzlX+VkJhvkLwavvwHdc7C0ADndcVRooLvOT83rK0au
zXEW34f8mWez1JAwReL0fvQ010xzBlYlgBYbkJLr/+IgFRo1n90cJGLJOJcR3CmVRI/8JQltJ4DT
j0zXbiLZT93AfhN161Tojil7ViuFWkR8tSfYOwu0phswDxyOiH9VNeXglL241wVaGu1Y3vmH4WLr
CDI1mlQ0tkgiukGKhpGmUXY21CFo564yq58ds6plCv42C5K4BlNmK47CxekhvfDnWEdoT150UKz/
QB+ERx+KArkmnT6ZD67ZQCaAYxDf9b4p0Werg9kOUz8cwWM1m6gBEr7f3XoYCV8V+yKDgM0gCy2r
ebD/szVZ5Ow9TbV938EGZZd2U99yr3TqQK53FhMR6XK2MnMAvkRgncnvVVzkNJidU9MiPrS+l4bo
gqe6a0gd+TD0w/WF900FvuBJo6nWiYlfTj6uzb7fP82FM+UUtuUqb+jZMFUL7ynOM6TnYuktxx3K
KkYiTtaPTtXh5pXPuUovjqHns6UyOrxX0gh4LosRnrul8DLM0eLuOmIKffnssDfQIBERWL7RsaRD
RqkhQeRUZVG5VXBwC9aKQaBvUe8qk/bIfkvqIo2WVQbMpjgpClrnhkacVQVQT73mbpyzO9GVeRb+
pes8w1zRFC6TWNN6v9WOqk5AvWvtIIHt11CZvhFlZynsUR7DJfBgwyz86VpysdG5CjnmTTgsU3it
Gm/L6hGzyAiEBFShMusz9G7a8bKpYEjDcoO6UX975aWsSoljGSBBBqb42UX215U6Z+aRDyNPUv0X
VIB9XvXsJUC9PU2/3syD0+3AYwYKm1l+7tOiGSz0xVeUEqx1yWF3MLgPfzhjTTatHZP6dV/tWTnQ
XHnnPLBRqLSjBXNeoKnPhoumFMC/yvup/w/pkQBkowvan9cza67JsO0bK5Q/XTumSEuiR/HTSHX8
enJ4VDGLLMM4upORjDhcw8NNM16QOSZbDP5axDc5Kit9h5IUPJQL5ZXtMUAkdeat1fypvspwjmVK
n3VN/kkz2/dCj5W+8ZbxdrxxB1XKHFSwehEeFKTXnymvMEFFPjOEXICJTPbBySB24Yi06f91CF5u
/CQVFinCQvR6Efoew9pFDiLy48KrWqQh4hFvXATgTsCqNYH0FHAIoqSQx0RRKZtinaDXAdQBuIQy
1PzZDvbgseYsU0zHXKmx18tEFw3n8WNu+qpHI0OlcyeOWR/aH30g4a+sRVRu6us0F/pJFPsGOCXJ
q0Ds+vejRLflOE3l4Gd2uehIDMuVzGb+mv+mt21tQRCNRSPVZonbTs/LIkEJnHWJmxbIYqCEOebd
wlP7BsTzg4vblt9AA4bLIWujZEkGqeFCXnwZKS18eQ1hbgQD33l9CQn+3tzdH7WQoPKgclxb7Fud
cZwwqvDjT47FbcmiapNV2RY6/9KIKYtAY2g7OUY7mDQZnQzGyugejSOcj30/AaP8MVaH4N/rhYY9
6IS6YuNLwVKfekMkeXoJ8NdU+NZsv/gDLPs8O8zAM24gPNSXqct5qYIe/4fGEZp4oYPu3Ue93TgE
pyzDIbKUsOR+MLqVFgt0fTXGgioWitqSSNWpzFvcWypZ5Wy+HNgHz5UAB2jQ8TnjLW/ZoUZAP/19
0Fydv1RZCzgIwi+Cps2lPKAVIxHE1HKBOcZb0TRy2khoDPpNgqMN9hpmW4kDsOsVdspP36yB9oXv
lVeu/ECXg17oZ4rl2NUvwysyt3DZjLxh2CewtPsHtWEWFkmv4qnf+elwNduCpmCJva1T+5cRcX5V
0l+45e9Oz4spBWbWhyUDWrHJZFtihfRq8SRwBV7btwzA6R165fwyHyE08LgqqVTrNlqjvLLVQoRu
H9Nor8YwjyGOgNIbOnQAxcI/Bu3fLcgmyojP2kiXmck2T40I8j1b5TwggGHxC5od3BVaaHWXotWc
o+JI/5ohdFk4rxI4kvzvKI8CbwXnV4PjScc0178ta3aNviQ7VDKAXMZH4hfKyVh6L8I6fNYUqruM
YzoQFgd+A8PVjf2OWeV2n42jNYRt55UbVZVnlMRJAjiJ2EJfekO4RheJT9GqoRxYT+6aB10J9Uit
HZU3T6GwzjzdhVVP4K2bR+5lvNmFg0KEQjE8Ojns6uf9SHGRpY4cALq8hVnoBRHNlRdLMUOmJ65f
a0jFRg1WGfOlcs9rcIj1I3pDOcN967tr/bpUxSdXiexz+uJ6auNVr/bXcXu5tB6eTBmEyL71mz6F
T+TI7HVc5oru3djGygtsvlb7NsFl2eGWXPMYHIcqPvFMP+qGPyf2Ip2TsLsnDPZIPU8XP7iEwmxI
rWECnoi1+YvK/ihLebeZX7sAWB8h9Piij3bJwL+iXjcg6thscH/v6Vr4SOyrb7ukewXdojzIhp05
UwBl2VHdKpo8cQc/FWZLHei7xNUy3UuSc0MjfEWzFsAw7/m1xeE5Z5u4pb9TkL07gyu3aWC5MUpm
xRQ3SIYXmWlXemXiIG+xlf0Y/YINpp4k2lmcWSQm8RFv1TlIFGLGs8JpOtp3Pd0EicstTjszCH56
E0iLd/bmwgl9cvZWlDWrx6qdF3DobK9ZowB8AenYW8Xoi1lg2gYQCdpEOVt3VbVhaVxvzvz0DwVH
EMt+S1sKo4s2OqCVh9pEQnIUsBh1QnlZ2kjJBm4hNJ2XDnB/Ru7nT1pdBymoD4y5uOH4jLyHPofC
7MB/K+X6gTlIF2PU5QiTTHvAKwwAnOOZLEKOll5zqBtTJE0mikNkaYBRyX6JebuiUrTaEXgL5vjg
rx3JpezTxNjWIHw3dzbKrXCx6CYe7m/jJtoPBi4NOzCdiLnf0zCExnc6obAr8PVBJ5p7YZepBb9n
e/9LX5jHJaCeXA5g75idrFVUqvYW8FtP/qLp1lOuu9UiGGb+BZDr6G4U043L1WoN3KNH492FmpMH
QaOQRh7oZCCqf/XF0roNDP+O3FhbsEyqh6oHiSnWeSZT1vLeDrWTypzQt2p/pHqfx+ta6pEEJqup
SqGympIZ59YGX5QYCLpFc1TBvmAwJnIfBdBVHkG9fbEo4dleUiGq8nYpo1cj8vUIAqrgaI0vuDqq
6iy7AI8h/eiSfZUOjhfrfdn0XyKLCvkLo7IXITuM65GC+QWlCdsEbt+2fgpCMRgBrDf/YEiVBWUs
zBjdu/5oIHuuoPRJwSHz7Ap8+ijA7lByo2gZHqHCNxBHbBRAKBLj5VfEzYwdn2LKuR8BVAuAWiyU
jRzzRMk2bcfirDcBjVNyFaZ2tFTO4HsGjtlYH5JzFIw2U0sPCpODZrnpPyCjM5JHUJ733CC6n97s
kHgq8z1xS5TiKHaQvSMeHAPZGgLVcyCvX07NnsHKB5qMsZradF0mqwz/JttER8+yC5RNBIL9oFsR
K9StDMSS/6W6laZqjMbg+CCgS60KkjT7SO2v1bZ+3jXPjhq4c4EJ7jzaTQ+073eg3m3SyaGqs209
dBCbdHhxRb/Mxge9dg/1JdAZI+cOe0JBlXIJnl/bxeNZLQ7hw8+YlCvxzcAy+sriK5X4jLD5B6HI
lX1kZUifCnt0SDrIpnL3zhjcxUdZ/vxpl2W0AgRrlGqqwc8pnJ7zVfbmtkJoIZL86IPE7VbseuGV
ZFLHfYTH5e/9Fh62UM/PMyJfy9Hw1Pn1h0CdQ5PlGN3EfSt/7bAfSzVVZ8n79Fc7caiNvi9YCqal
oxksd+5S9Ra4TlVb88VdG+4KI3+BpQxleXEw/x8QCzORncU6eTqHpnIiFHdJoNJK2fOBmgZZgrzt
Qmtey/hqn0R5onc5AaK2+rrzmzpTBPTlyoMM+xxQ5reVhQNi6tj6BFcl4JPN8CRSFswZRMN/f+T0
MXLIaKMFFEaJ0X8dzuM1G1RkOfjo4CLRUJojxzSfalvyfV7xuU5PhBS80yukeOvakothdRmBrAts
6wlRonMOzjAS9zLD3HoD+dNC79IFGqjTRDgYZvGtmoVYTQHMGCCqI4loRHHUEIkqbBTLvUfYZ09t
8/+duiHvJQiPd5OtPJJIOPnQJCVKtuWYp9ADep/NwokfsK4T9Ive7R+KK46QCxzk0E7Tcsvq7/Iy
pKeux32rjrUA/X7CHlOjLmt8KeBAxqlpDDydjPvGmOe0c3yQC6m8XRvD2s7E3/Cv88lf/Yfn9SHI
qnt9GVTADoYGWlQGKumKy2pqJGbWwUFEL/gDXBocuw3c9P1Akn0RpyEc2qcPtsrdIEewXA2eVAFP
W/sX4ImuhmnKjWy5z69sjwyts/AIqzNbLitHuMJ3wX/0obpTb3pz+Jf+KZbnPoMctfQw+sYbDLul
emjFFwJZjUsNwGDCYUgo1wGo4dYrIBEVPrkvcu/9rZeR7AfQ+NEnP2WdDrO4w4NKzSHBT+f2ViSQ
/1sHQXy1URlvpQHb1yO6TXDOk6De6hzoghowANKuhL5QxkdgE9nOxp1fmAwLzqyiMkZYDLl+Wg30
DlEvB08ChQtHmFRHJhZA8H6ryLuQBTbXyvtPKvEiM7BxMbjWlnpL68AbRH5TcJxsVxNZ0xyXppT6
njvIqt37UaoDPlrhUGtVoQptxSkgBKZN3JwBuHnYcxxxlhn+eAZf/Sa/Z0gPfG/DDNsjRgalto7J
b/HGp+MXoGlLpkFLzwaX7Q4R6T+gFBjZUyM1MeTK3GX+PUFiMN9rUfiQ3x/YGBZIzGrzHvOFP/ek
FK2ACLxPiTZR/eUpZ/vNdEfXGYaat08wdin07P1vIwZJQWUEz5XeGGhWUmWcRR4zPGzgiy4csVuD
EafkgnpDnkJiBjATJ70NXdwoisuvMPsrRfhLCvXyHLUuryyrJKyb+0SWpk5EslAljRhA5ZsX7Opg
CLjxjblmKhYtNcL6zb8vAZE8N9LysjjUTajrS7vKpMs6giN5sWyt+W7YvlT/iBSMVGR8zZbWn6Eb
FK7TY2JINAChwBqpxy9fLzwC/L+kh3YRhJR0qtxa4Q5lgn3zbqBFiIeZyHhlWnUkAP6EUvlILtX+
rYJJek9BxEI4qBKGm6el/PJyPaoAblARaGhBxUDfxMcfDf6evU8eprdPbmyr7Mv8CGYPCkcmaR4g
7E5NatOn4hPa5vZpwyzRL0r11Ur+EczfaiNlPFqw98c1P/hjXGwp7rf5TJVvQXQPnhvKjIvYSS8x
P4VbEMi8gH/NWuoUmPzdvkiRzP0YPobH1bxTiA0F7whY0bQYU3oKSQ4CZJ3gu3pde/FMFfqtn+gi
WdAtAkDbNB+EEjf5ak1NWGAibXq0i6m0S4XGFJx8+552fdDAeDft3a06+P6ddgyHSbPb6GSFXjnl
/s4xrUwcpLPT1IgJytoxU3x29aQiiSr7vE28KWSTWhKn4q99lwBbwpzn0S0rpVFgw/5xXFlMPOPc
76tprXBrzr4apnCTRabo4f1Cc9nyQfNxE0e7+4ZjSAmGFBXQKRpbH/Kbu7EnxVcZmaW7wCm6wJum
9NouaKh/20yzBLpH7x3/ZbzESegxPrMxn0Hu8fY1+qSWNXDNgRBGPlPHetPPIMSZbkU8Uygi6Iy8
GHZyK9Rbl5h+SqQ9VwNI60AYyBh7dLTsYaO4eBxrTrCuztqMDC+zvw3VTWwW3eoyp9KFKaWkOm/P
YrMb++H0aOPnt8KHLwFxtH7EfUbeRjQCp1Cv4XzUcwBQ4wsW6+llG5/CqU30N9McBl3bt7/IqQu9
M/e/Kz78On1mQTSXim+Jq6niq3C24VfNidu08AwvcN2dgRR/59rfo/2uEmnmq1o5HRU93HhkYZsM
MkwpU9DW8UvBi94CYEcka0hmL1YjYB92rSJGnDlap4P+OAPOcXfw5K9pPc10UUckyxX842DH/Uje
umvQa1PqdvbXJ62fTGZZ8Ufgbw+0llOJsRJ11iy82eGXxpOxwt7b46sBL6MWBjx4Objqf+0gAJup
zW+Y91MwVgI3r+ibAEsJD55AiR/ZkPmO4gD+1tqmRNEs2+oCts6pd/mhk4YhHoTZFiMyEx0Dju5A
sFsQlkmK4yLLmTBvoDlWjAr10niuGwk6oh3Vnwo3xn/NtY+UsaE2kXkQD7b3pGqmemYxGCeC1zjG
PZM40/H28N1VVtYN9/Jr9sS64OYjD1NarImR9aaznekDqdTlxVpPZIk0WsHRAXpD87mGyHG4CXDM
NQqtCdhimqJpqUInz27DHtCMoEDGMeDaq8jenBnAzrQb8LrawKsNi42vedluus36YNEI5nenvWLD
Cx+MqgVhTfPb1ov0Q4/mmQ3KYGfLkF39jlfG7FRzlwRAedfr+Oy7HxA5Wt7lMdKIZ5bkUfF3ELST
UiNzxWaIxBzZbm4bOU4jj0xk0gwVJxRfVu5hZPsGKaNF4H39PynytLVjgT3V0SSuFSWNwaELzgeg
ft16VCB+9o9zL7qhtNHtQdqNFjGKuWOmvXYFzfTebbrNtiWOXBs5MaeBtXL1x8UiuU1YcTRFMaj3
ygjr3bdsQTKQmUlmemzw1OS5aLIStMWYTI6oZPEHHmB5QTfBtXQJddbvlGuxSp54ANz3D5WzMTLU
1+/Ou9t7Q91PPFQhbkDH5Sywj1dwC2MB+MGgentL5dlfRa2PfH9wpVIDJzKm2qUuiz7lf5Cm2FwG
RQLvcQZIwm3lovGLlgyIf7yeHq/iLKtnhl06/2UtL3aHncaMFZrKp6tBBtVM6d2WxJl3aJxzBPEp
4lth/luMS9Q5AvEYWk+J63b3AOMYYvKiwzESAPeXclADSK8w9Ds71aqocfrCt0vrd2ZsyaBrboHS
hgyDihWltRF1ZoPpeJ5vPSaP9kb7Y4NBKmXgoJbVOkD3eV/an1cNc2WADRNAG0mKtGd5jZqP7XkR
rKvZSz2QEaBxTQ89fgdLkiMMTGGB+XzPhHajks9EgHFbFkQi+RbPKS6SfGg3hFPNzNw/tE/iTz3x
ZZbmUSZgBDVfWWmChcbyCproQRGDOlL8ZGZ7U9mGpTHRR4YhkT/SWSZmUw9z959dLzY2YPWyCm0L
arSzeFplb5rBmbpOlWYyHyl+JEd82j5vJxBExTOrNJSmjKsIYYcctOB+F4pDbOSvg1YYQltNJRYY
HXaZ/Kxv5/3ziCpPicQgK2l+9/ANoPma20UpbqXrdyAdA6exklxUq69vm5li7GOH/SSVvfJ+sJ8z
VKn0E6MbmmRe8i0aKk4SV+Wb3ugb9EVLtCb+394EWmIclIwJfh/JQls1/Dqzt52ztQiQKbQZtyvB
ZqQmywMkthsHkKqeXTlMliYUOWOMrFxSx6sXek4AyI+YsVYx2xDycFBjgBZTumflgkKAfsZQuid7
7U8bhW+SVlzuMrvDJxmVkyD/f5w3pkMrw4xRK17UIEGugJWjmCcVZxpqRu0PIphS3x7MhDWp7s5f
XD+2lfSregTrB07Fm7894/bNngl7VfrJQ8dS1m/ewDXu2lvAmw0G1sjS15l4ZpvuN9TDcpBFVKnA
Cz+91qM8DWMuE9Ay1ZrJo4ZJXD2t2c5DpXbgCqEdamviSXFmbqsorIxTESG1S0gR6kRHO0WYliJx
GJ2npoB/7NiLsWG4HiZsOLkRRaYpf9sGwnNnLM+tBsfSauT+ZKDUDRJmYXyUwB8uLT7XGXAFcz5U
U/dE2iqjs7SYf4PBEkYWdRbfnUwOWivZKBUkWyTMCcSQA6NW7MxMLb4VUxUzSB1VNGdjlxfzU1BK
AHUI41Sxt4rdsH2zfU2aU6r2L53Fw4POED9AfVJX1KYh/xrEoUPMD/z87VQt3rlVBNnG1Dlv7qxY
TzUROPMxLuoUyNZ+R6sXxShqbDpwwp7A2y9/p+vbvjoaJZpkCwMy3MP+OUEXq+yGQjQxS0GLMr6t
gUBv3a2BfcjuTNnjgNr5a8dKxmc9tuh323jfYut8cLlXVfSqydQaXUCa81h5uQqIpDhC3zsxEXed
uNk8qluOBx/sZjO3EzZFnNT6zN7I5AmfeAtC148AeMQ/snWXfiqZwL7ySeY1RmginvTN7Y/4MMGd
nZvyUee5KOgqPBbOxkqXcEi8JD22JORS1K2QydTLaaNQP6eyvryhyObvTYZ93jTY1fuiz9LlFNfW
z7BGxBLgPY1wFYkU0IkGs+ssi+JliDUkJhl7CC7rLngR8eaFIAzkD1S5bgGJbtwE0mHQwxjczgRV
XIpip9Vi2xpmnBaF07E7txUG9chD2jbB+6o+GgKH85oSjZucaAOdiCDXh8eUIPSM2p4UDRzt+3qV
8yObipBaDiaVuwOagsvlH5BUjkWFaFJjTi4a1jTtUuNV4JlvlcbSGmX5pK03ZsZ/F4nsee+CUYl9
U5vuDVrJKmQt8H3tif5dcwWZd3XRyqaZ/v4OB2hqXUcKLyf0hF1PQYMFTTQo32QGvvqi/+ftJxsV
YC6+mM3kbJuNf1H6gT+zRb/ruxg8PLyAaC8XZzgAJqdW+c8UrqFbIDHncNaN4uwo55uBqj1nJ4iG
fzaJ+ANHtCM5o3gLsIFqfNJlNaiefm0YFvDv7ZDPpetCzuFVdR/Yh6OEWjeEsb0H5TOeSjkn8HdM
C2bpbEmowfCXV1LdHMGam+kEAvnv4lNz88k1UEBLLIU+LhrgVM3LwEN1NI6HMmlAMT3yAmPhukNW
IjihYUkHAEbynaw91ok/UdcGq662x4pVL8F0jjdnCuQEjFjDjV3aCCWmRciZI2nTGtr4StYSOuSx
6zaJCYoy2c7EzdeKPbgrW1fOmVGhzgOlhiC8S1h0bCVHL3iTf9lXbWsdd9qsbzqVd/tD1TirjBSM
f4lRm6cUD1p8KFJS7KRvibAbz/u/hWhvgKwFMzQzx90Qww6qtSxRxCAJ++Ijg0AqZbL5dWoNT7AM
8HHi5j5hxrsFrykSHCmRlb+hTblT5GYTmyfLQrPaFwQbpo3ddiSgRd4v4kKuKwQyuzSy6tDKklTO
Te5EoMG5WW83qKjdOgSrb1ACzqEtKFT0+JE/r6RTEwf+5XgH2vRNReC53mUCQ+PvNrqBvLbpjkPQ
K/nqN9BohaC+2fqPAhw3QcqnKG4xXiNQwJd80W/xBUOT0oKeTNPkgEO/rjnCKmsfxQSruqe81XId
HuYHl8B6mD0jXxZ/B0A7jLo00j81f1WRvrMv5Ej641S27ljBOOTAKvfbZeQ/FpMo6SEjjvwDPdTr
4pDJ7c8fI7AjpkJ8wSSntAWEvdsWU2bDpb0bzwa3clQ+XM13k4z+ge7sTAMxY2Z50J4ulNVmOeEj
cxgMrGBR8Pr7MAIwcIMNHupJNoISF4Qy3zpBYsAcq7snm5CRpkx//1/xhV5aF3SnW6Ef+BrULtYy
gaINjrmUGGSthvjj7ct7BGRFeY6qIQrMycGr37zBsBBGY4Scqgnj5hVmK9b7sedNmeF2nNLRfFvg
oPl4KAN+CTxOvbelZjdVfqhkvjcIvOu8ql+aiZnY20sDQV2vIqxTF5m9d3Dl8PNYakv42drdYF9p
VUovBFsWSvjB649EClxHkX1sFcssn79TJf+MJ0TPiFQuODjub/XCOQtsj7TXvvHEEGqUJLXRKgyi
lAddY5WY9gk6dTXECgTZh3vYb4csTl3VIFdpM+cPc2XSdGyubEULQe19MzIjJ4DsIm9S5sY+X1k1
S1IQ6vW7tm9GScqf8v+PVOnX1/FrSEfTkCYKt8hqUeDGi4F7uNYjtCAphGwILnvgaDlY2KOFcnFn
XEButIebKqiiLb4qkLdr/E/Xy1cNPWYAiGDx7mMBmvJUWGSRcCs4sJn/qiR5UeM/pwYeLpo/EcVJ
cp5Zvr/bST5EoqXvHYCQQAAcbH/6fAJ1tRn3gvUoesD0WK1FDqjk3e7l6MrBKOX4b5RPemly9IwG
z+l8uNzqf1nvmisRfb2CwjC3Ec9D2lADn/b+oK9kZPfLHqhihYd+R3nvMKQIxkGEBiJXMRRhqo5V
rkB98RHQOSJTYXMqGdTZ7Brqmgyu3PX7uEZO+MJXyejnoJQ2vUwMW1n04OUdMqBcXnOB3lqrbpLu
F45rQz981EYqqIZWT9vbXmamW8DThbV1HcBUNqB+JCisolPZ26dAwqhZJcY1vWt+ddfdtTYQMUQZ
3rXWSAOUlw8w7VpAOPkn9pE+ryVIWdGfO4Kl47EkW1ods0GONP8XK3g7B2aEoydiQshF1AsrZMaN
LgZbR338uStI7MJL9qLWkdIwHrYml6AqlZD5DugCX6+HytBHHAU4oCL1zTelmvygTgTi5gPJo6Gl
zIQZaDNzBEoSYFIFvGKXe6LMU81v8dXN72p9qechER+u5FsMTZmHK8HaptmXGqEjjn3eFM9UtRN7
NrX00nyAATQdFN09IHzXqoNNT35j3LiWdtDz7oVsp0D1qn+hrzdPh7B4gxODtsDaDtPZVSkhbYGb
+oOrn5oQC04XIP4nM4RpbYkINHKgIW9OmI/O6mKTP2tOr7w2ZvmcLShy9AsE02qavw1chSbyOe/L
b3YlTjsiB0cecE7KdbCJvWFKx7DAnUlBJ4ATOaAdaz3eWDjFAq0KAp1au3TXt054UfMGMwmSVHqM
Nvo1IlmUkbwYJ4x8BmIL4C7CrbsTNPrk+o9aMp7hMCMmux6EIn0VioO0IwNHaQY4q6R62cuNQtLM
fI/Z3m9VT1K2u4gQMWnNDMvAPoHmFv0dne5CSRECdOwNbaPKS+++TuACxNaVUmrxi2bwENGnuvMm
BAozVLNLdKNaeh/LSit+uY0besnJ9PnpzqbaX5RiDkId2yjvk2T4y14ae2kqGc6c7M160Eiu+N3Z
+tdYlyqHnv5cwLME0NSPtFNL8gsfPlWj0/7PerTk/iPjHe3hFREVWpXb0vomyXLjU4To6O3qS82p
a1UGBN0j6wsr0kfyPaDk5Xv4vdSRJ3QF+AvX4Z2OTAMOZX/HEDws3jJmYBEj4EECLKxAygl/eTSV
Ol1eqhCCR5yX829k13ouMzDLxdcbeY6yRIacpiH7QK9H9fccYkVnu9IqjMXXzDI1JU0LT3ArMRUV
06mn5J3M5f75wT88PD3RIjTTscP4ERvmhR/Ul7i243VpJQtGhdXQxB8cR7AfTUdCHtevs4WGpF2z
Cjbq0wQN3aZSKRTtaphLI0of4ZKSgyI8ee+L8jUhPbF00e2Pn8ZeYqdJ/JTEa1hRJzR82/8Dyh3F
vwgIfGvCsGMx2FFtkmI6rj+TUZjiXdXs/vDwAi09uU3diRD7GnAR9TPqovPebJvuV7QkSuOSOGrl
JPGr/Hnvoh2TCLNMVrgBp4cNttWvMYxnfpLsqUfrXRzwXzuMLpI7lsTwESEkSfvnkKuyy/hewKRS
d2mJ2msL1YNLFG8r8MQaSrPh6r5oyo5Iywamx9okcV9ar59Ko1E0t/Uj2FHV1wsbwOmRrrhkWxuc
rZCx3iChdIIRSG8mSAi7aAnQVdlx1BhVcOIZ/dl+gALAkGtg13bGrwjUushymXOJR2gOzl38n3nl
rNQaI15lI+gRmYWWpKoiKKDyJpP54AY5zv7L12ZnSXxsoyBWCsx1kCsOFUy1ZIx0qsGogjmWuCLP
2JMAWk29sm3sTDjPpSNsQ3EZ2Cicc20Z99OlzWtHZMnyFPIc2RmoA0eu0tiJSFbm6qps3wU277s2
uDsNGsHVREDiWmR76yQU5NCXKnCgyZjJsdzQLzY/0VwgF3dypuDuoHLKt5DRPF3y8hHdmtKmAwRm
TUvJjjiPHewoWFtIUltfBbbgBjr/MUwA504x/cTZJMI4LFiCYYLOJdO1hGzL7G5NQHEJ4w+5YUAl
zJ5q54ak7rv9P52l257fCorsvGPV8pv4iVot30Fr5JmfHF22twO257iR75YiYlEATzNrZ1oScBA5
wolWKzTTKPrUeTG1Rjq8nyeoAsr2fhEWzMmYSPctxb1lLZsWNsfzTcRYRC0DS2/NmHWsaq3vC7O9
0VBuVR+VE/W0M2m2pWDJlL/cwj75zkrJaQVYPs7r2lyTYxnQnxbSwJ94M004sbqk6/pmLrQKsZo3
zj75bZgCZ7dfoMtsWEP+43p4on/OIMoAZGK3IYtbUY+J7QZPocp32YJdHGzMvGNEnAeaSSQC68Kc
/bXoPnS19kdFYdBQqSVyCjVd1Zuf6BT0Mbjb2H/Mp3eerqhjkKBNvUN2wu3v7/CJ5vWQt+rohtU1
j3A3Cs1r0n4l/KcBJqnzIjsETTfKkPp23p3ittwVz+fr0gANAiEoWiufJsEbMZoFsPtxmqGZUqYW
9CbG59fU4v4nis607ISGWONYuI8qsUfXGfYrEl6/21tjYdkq8lwAAbkNQOgk0mcNoFN9ccxfbmtc
1kuqssnHTpnR+pkLA/+FWXJHVeDe6W4ZHcFbRhK3ErJd33V4VbAsbPONotUtOPYZC6Tl9fO/EE/0
C48iuKHUr9DKRQtjPaChm6yBS96TEaogZBPdJ5G2wH2PUxAJy4Fj2XLjHLXbZLRJTz3cwWXRGJFh
AjaWmcxYvnQhxwVro4+/Lo1PU38ZLtRcX4X8xCdLrwSs+cFF4HnuLvt3qs9MZLOFQn7DvQxGCa28
pRIoLGqArz7uayUOoplYSQjlkP9YZ3LigmdNc8q45ORzrzz2lK0Rq/0kfFCrXieQpE+RDgqVw8sy
nAq9x/aXiyEdf4fhT2u9xBBvwE3DHq0pfmrSJi7ji9MGEhC+Dzx44rJZBVvqX+IZCC/k5WmiTuoQ
7BZQ6StkAmuxWFx4W+iPtDSx5tSqgyVAZdeW+Y//gH+fIu0Pt/AtrM45c39jeG12S0GRqj5zr36K
UJQ03JCeJoUVxHc7y4pbN6i1DE5UFj2O/BzGHJXfdSlzPBGv+X5Jq3rSYcvzZpf8M7e0m11bNcXG
0sde0fzPXf12DMnWIG5l2bRlheRqCPY4adL5mHs+mm0PFqT2TkgDESn/v8USuWJDXszUuq38ntb1
8qFkpNKk1hD3cYWOI3W1X5pmI+8HbpR0NJ+5lVf+g8WDLRmu3wsYcszgCb/4X44M4TTIsQaDpuoR
fz/q6B7rePM3CfxAoZFE3sJn6GyQYUnNWNlI2WQbi5Csb//0keDp6NClMoLoaW/MA5dqTcfu29Mc
Nj2g0JZWQhMkSeo05ivO2SAX1FiFpzoe9V6dEfCiLrn6898tcGgz2v1dusupe+IqNqR8LvvJ37eb
PTYK3jkJX7yBMB+8tG8fUNUXEGmT8EDeME8MQMTiIklui7f/v0TKlRSNjuydAn5FzjrBqzfqL+Mx
3sSgpjKbDXqz1gg66hcBck0qKmakBUTGFCCyE1nWh1oZM/KAojcgg5qIjE56B0YkLRhNER3vlgSr
MlER+wQDMjzZRfqwn+87xZPXkUw1Mbu4C7aAOyvP75IHOe8vg8srtTdP7BcgQLse0cw/1cedsiqN
xg7+AfqTdpXv+ztwnEb4e3UE6Cvm+PgScLCUCqzMBrB9LQ8FBf7K5IWZFKhqHpvPNUBhKQLdIiJ+
p3zi61yGH/0nRDYW9uBOzbHHoMAPZKRqnR6lE31pObGr4/G+M6YwZwl1K9LAu3pFRDX6iL/JsBAN
n81CFg3Cru0mWzUFyJUuG+mOchHEaqn0M8X6144cdeTPhudtt8ReGUFTmdAt9zzpRNMkmBvGPoPq
v2gvV7inGn4bH7MgDPw5aG4JhgoBxfbz6KXRHk2MoT89aYedI6e8qwOhmTRZgHIfT0RC3Sxg00sd
42VFwgdQCKGUE2udhajTJTJNa6RrQK9vnn2QNQFhHYc1jva/RitOD+oKYy0su9uAlImeJbzehgHD
5Rql5yZpCe396Nng/NaU3FE9U7j5Wm+vpIo0xgKp31aK7uL4SisieMAtY7eT2vd58jNrctt7Adw9
3dlbtAWB7s6Sn4iLtIfK36vwHqPljnvy8WskHD6okhl/lcIJMrtPQiidFtDWuR/dAC+Gh6soCh38
MD1YL477zv4m9HM+SEm2hKF43ZWC1JcoY66IMtKaelC2q/7RfAajLNT95C/Dieg/VtVM7P/CdiEH
Yzs/zB8t4+aIEpzdSkBTd9+KBC5ADpyypXR3pIIVYJ4BLnJa1fzIawwxL4s5wBukiAJpGavMNRrg
yZmdGuhoDTuvI5MF9kZXf7V4llgcYgxCV+klPkrovJNtKEdYpsKqTRgRHrWgGEKNtqFnZu8yfEFz
rqlUcl5lCscAQbbvi69+woVau3ZZKOZxT0UA1XgJKjAja48tI17X1DML1nGBuYd79MtcbZttUv5j
BApL0CMLTBdO/cNgh1+AJJj6RHytCZdLoEzlo5A7TiUw+XZ9xP66TA3YFEKzmRrPheduyzVqcE2Y
ajDjLVL+2Jvc4KQQrQGeBE0vWuOZbJhM6sPKJTc1EA9GUcYk8XI37p2AvNtdd5VXS+90zff4pAGG
qy1pv8OR61RaJxzROPqA71bv1revhvHhYqUvvStMwun4mREf3fOwArkzh7RSL201cfvxACabbhJ/
ZZWRvNTfL6vLeWj7opdAKFbea0zyO/cOFAvPqm2cPvbIlJ7cITO4saemZofYY3v7leMc0tf6HsmE
qgMc3ZT9JPo6C/9D08gNXjiaWflIIxEEBBQ7Jmvtp2HmWR7Y5bt8dh/G8D2PM3YVz9Ew5cYEVTAh
4voXvnJCNZlFG/ED+fxhRqYrN2muPxPcGMRJvnkWGHGk97Ew0oXo0RBCyYAn+esE2syugXcH2Br2
iAn7YzPMbuUvTU5cnW9FAb21nNjvUAKlZxNB7JZEORSXOmY1zAcDEEhRoClgCU0KDhZKnjIhuLV/
PXI0RHz0rzIYKJ2jAnb3wjpQ6YeD67EfOozH+y1tWJz84nFcpJwLqlqsBA0wdpQyRJuRYWjeefAY
cw0nYVhqFJrbPZ+VJTobw6HHjjhvP5oUzEwUiK/FBaYT5yUzzg6+Idw7nO8SvYRVf7gts5Le/jGZ
zclVhsXJ0FprFT48nRidw+fD0wNMAGEACeVf2s0iPomeou+SW0Ly+dT0qFLfVANelCxrGEqe1YfS
jQY9MBUdoQ6MV5N6ahAWNyLbvVdXMZtkyF/1FpoMn9H/5SWnMAebBsf7mS/ULJCIikdt/HZH1kJ2
AcA5JKoRDP0vQfJ/2lIqm9acWSw93Q/js/tqbGkclgh5bkDoMAfeLzUfMbRyjA1zXGxZZctlYezw
1Jmj0CW40UM6yRHYouIbm+70MkegWjT/LNTPKX9MR8SA6dK+OIGnYVnXuwCrdLMEqpBEkpqg6/Dq
0YvcsRSyjBp5Ri2GB6JecG/6BNMBRp9kD5F/qf3mQ/3RjZwkbknMtv1EDDLzA9OKmu+plbEhDCpS
iHoC0Rqs2TMpVetKfDZie82/tu+dVF9H9bdgH/Qam8sD4Skw5Mn/QXiqLfYO+kfQ5uuHavqHhj35
AbPFBvK64uyICghjJ4nwE3mCKSdn0/9XiVSQbDJpF2fBCFiFqOV2nUhDwWBnSzbXWxpGATx0bHfN
CH+mnjueIeHm92vcZVxE5Xr0gyp/2BBiBn+Rda4D9Dyrj+XrT4N0qLf3c8fPVTOahcgOQBSXoyVW
mnSqUcNNeEtnuZOvecPL3BtWvdLgFxS7LItbzqe91l1nIcL0W6VFXt/y+0YXw4Ev5GzQXuOLg/SS
mted1LYht/f2gG/XgH2TDG2pu+4/X+3Q4l2JRZDlzmkCjJdSBLMJMNmaKlNzUOc3JCJOyDRH/3U4
zhxxtHEbbYnuzv9gss8wM/pFMf3scl85g7/Zg4MlGJbDi1FrDY/F2XbMKupxlw4B9s2q2GwnPSGM
DwA5c46rJWGy0M+BVLToVgOMKenrCxchc8B8igt5e1gWkmGiyQDMXWSeCd/lzJpVq5hAS1m6m249
Stikwd08tqZw+s75dswtKnG0HiHdjzgqjClLu5H4pcjkbPgIVETHTY1e4EiFn+5cjv5aM2ZfOpi0
2+ZuYcHnu7s6TY1CJN+7iEfdAQ3XC6Effg/wHHB0WXw72Fx0838G/rKFRH8ufTpJjT0SJUwfAOem
vKCTwSzuMFTMsfFIoQ5Thj3FuUyayzDchqZ22iCTJebQryMhMESjxh/FO2ivZDyJwc7p4gwvQ5eG
ybnIvah+ipamhmhejhnN/69nufHthNyzbPXc+c9scynZLeemdUpoisNj1H92wj7r+wBJuhvTNx9B
nYAywHJSc27FXqxeMkZCmFSu+dGIP9XzOGCfene0tBZ2nKC9dBIfAhn/GnHi3q1z1otVVBOhFGo7
EFzSuPHT/S1SyrVDpQohasN5Iy+Uf8R+6vu7pD2cswkK1UI/vyclLehXamLQE9cJIXRvccsWI8+h
+5bwD/yQFTSYrhyDMiaW9wbDbR1/OZerDQNqTQUaAIvdgaJjoBo6/CdJGTuP+sYPlAuER8XNais4
2qnbOAFvXl5OSXS+skaIkZ0Hdkt//pSsW/vhajG87rBx+chikRBLQK0wiBQwyTO32x4ZVVk5owKV
ezcvS6MptBTpAW5wGQrSv7ozAlSVgb5Z7H3mrndGYa6qiMloaG99B62KbqiqW9g6mcgsfpfPkAqA
+DWbEAyZEz7CNTwzPwUhxU0/xdSJt/Yqgtt5aEKYdicKpJEbjQVO8r1Fy4LDs4xLP+3+k+WKIUOx
OSa4Q9mXS2N9KAcL6VDEt3siGNC7LKSSG71IIbyTPZu6dV9YYNlSxh16NZTR1948O1RshayuJwLI
ZOk7ksG0FJ0mCR7TMRBcpnIE3/c/FWmsd2ZEBar2uqb6LdvD+OKzNnpXukh4EYb5z03bAInbgmiu
OflmB0Sqzp78jzU1OLujo4Gx6htxmPJ7DkeVeDD8xUPhOP14j9SdpqEGh6hkN4ggn1/iR1eaUr6D
NpYz/4QJKQABElxXCnsKoak/NW8+i5bYZqrw3/j+S8DCd4crnPGA6L1LQXVq6z5nR4MnVK53vAA5
OLVqzxYgGcmWw0qPdluMrTB+80YuQoCG/qnicByV8ag0Q9SxF0hbL9HwBQTaSVVt2dt3B8GYdj3U
XKHJsULuRwTPxB1xsvNOeKBupEuRJOeg2rsCqIioJ8ww0djkZfOAu6+9nHLi+BWjqywlKzxcI6U8
qRYt6DUT1FJvuSrSUeHQJMo8zVbPPmpTLGfLhbp86xG8r7M819XBdw5uQ8KKJaXfr47qekdWd8uG
BOPVRNtYxeRZUxKJ7xucp1QaoT5isqs6OjKhCHYqZDJGEWdZZ9zXMmpR67r2k/L9wWgZh5FmkuiH
eGthuCOSbKXZejvzd9eqv1DB/FXYJNHXEUcQbXeEpSS1mSIi5Tf9Yv6+//tyfIKbwSyYdnMYP3RL
it8WQrwm0gslJRFMpdsh36qiwbdX6vGRXvFzLfVCxOIydPkN/mxtkmNE/h+s9x/oe6yUw3YK3Jh4
3bhcp1weUn/XM4AY/ebgmkkWWJ6SvXgFxoGSDwjHmUQnt7cA/C6r7f9uNdgIIpmveqjw993YsNQX
rBiaoVvccHBB1s2oAVj1csNq2qYZyhqMm+HdbHoywP64sJjjNzUrCnrUyy8Sm/xtLs2VU0sa5mKq
wrvI9id3g0DuG25wiPgg+MnzGcfOMerCORRjaWTazQQDs671XIf/T/RbIGwFOP4/OHqvAqTo6SSB
Wz1pND4rQaA4f5EwAI/0vUhpUrqxjn7P9W0WcWTL9uKMyYqT+fyOlcNHL8rcraZ3+t7b4FSR673x
9u35RWzhBBRYVnE9r1bUPw7yvb4iwUd3bIhAcSzLZW91AbWkVVXEKqTe+XGEIfUvcrK7p0LG5wSQ
06ga4ON+rQloLhnOsbWHmFis67Kscww9ikU96dRLesbiFzqXQtq2hwtG/d2vOvL1oIDZWSvUkd87
q5P50avuUoSEXDaDGDu5bsABJgGQjfNp5IR/PQGv1jp3uc1Fo5VRDKuc2RGsfJ7Nb1rrxu6naqGX
bVVMkBenuKy/CPlcf0z1xDbSHVzM/0HWpxm5U8bmNAiSD1j9yGmhGXM27k3m3wZCbrG6mhO0TdCs
B5IADYBLROzw/wX7ycTsUl0n7mt1g3so3In52Id1qLyOY0w1CA+/hzp0yodRj19GgOyeMjU9IX9j
gCARz+UGR5DtWnWIS5BGTK/gx88vsiWS7YZin+wyjbxNrO37V8BT4jUFk95GFAGw60f1xYJYLg0I
km/n7rv+sq65XHTQWbbrqnXgGbKSL0uowgPLcLFhSZVKBkaZZ4mMJgbfHr0mr9BxR/FvfN6UE7yQ
N0ts30MEiO6MUuIGDDugvrXUk45OjvTvAoZzoQ/YhTxhIfyoVVg9GaJ9uD4AuQhxF531bugPlJMh
g/NJVIthAC3kylJNW+HDiNfgpjXdhMMK0PUKrWZyXNgtJUKuZf/Y1tig3w1BMtO7JU00XGRhnyli
a5HycWkF+hEVmR7SebCNJWHmX7ERM/dChKJlLtmT9i6M5zeECr5p36T8iXGcE0y+irBpJ8/9XiEe
Cmnjgzm1QtsvxcNjNZSFC6PMErSBznfWsrrpDSViVZtZObxb8jIodTczEC71vY+kd2WE2wLb+Ho3
ylkNQUPQZnlmTmIiA9rAWG0pLawt+S3oaKXRx21PoVix6TRa0FsWsEkPgZ/LwPe+dzhIRKJ6EU/F
8V8EDmB3qPz9rFVbVISAuVlNjROQsdcAMdF5eAIx9nVX/sFOb6WNLtjy3Qdvoenc4tjcH7uvgOGH
UFARyPVMGQ9n4UzbW8HcXb1y/lptcbgYOWoqox1CNkn4nbyIhqKqf9iIVBTMp5iU/neIJlgIlGd6
j19EM6B0UaYHe8LtxgaElu14+cRF4evg+V40bgrABPI6A5T83n/7aSuT75k0WebtX/WJ+FYGLklZ
eeMlHyEaxqNZF3pfSx9UGlg07rZf0z+wIwxLEcrW7cDjgQH+88+zwlfwV5rZb98D08XOpiJThKqD
R0GYW6i1GqC2T2ILMmmnjR4A1OPnlSqjRmpAhrmtTLld580K0lm8Zp3QQP5j6GhqPYkPgu5CG4Gk
bosXJnZQk1caP33fvZo/3tT+eHDqHH8vXl9CmDmkL9NCIkF2LU5EOAp6F5TWZCg8QihfnVcx4upY
QBScc+1f3j2LKs9j5eQEgzIgLRmo2VlO6xe29PiIPtiYT14p7L41yVIKnUlQRjzOwjf8L4luiWXM
EJdu58G/029NXWn6qDificgU8/61ABUgxoUBm4BLi5scRnmuMuZqhF3VukUB0QL6VfxI5+4ilpFW
6T3lfi+E65aF/uMrKMdHgb5zhHn0aemk7gm1RKOitJesBg29+Ad0WAkqWQALtBD7FCe70JZ5n0Op
FGgagDsK4+LvbuLeW8Pcqc8nysN0ED4Sa/GzTkg8Px75SEHG8DpW5gVsHSMbUjuQM167sSe8M98s
PmRiTKH2rd053L1tT537qGCf68fYG1isqudQhUqI29nsUCmnpxgYIr266jeIecBGe2PeLVErMV0Y
FH4OuM/TsUNKDLaZb8MARw6b0+AaNXkHjllBf4Vs/Euvs5doU64X2QzqfMn8VCofx7ekkBEbqf3j
p8VcTNdUv+I1ValMBdKZ9Z1GHxGZZqfYynk4ZNZBXrgGBYiM1vv39asUe3kiIOr2yf5RUQnU0lt5
EgIMO6cpmQ8MMSZmvroV7WeIp+UK5BaQFc6GPIYrJk0fKcGmBjKLWo1/4MMTFyvsocUMRPnNub5E
dxJs32V3fi0gUi0U/EljYm1MSNsVLiRW79qQFftfz44ep232opgLOC3P7l+DIuoYzF8q4NOn1+cu
VH22Pd9kZvOKjYfNEWNVmOTtXClLohGbN+0iJtUknpTDGyqnlVECJShA0tgTXRfaGZnrHzsUx5R/
pYT5++yoasrIqUyuA4J1O6j0u6rQYNzBqFJX+ii3xiIZbRNlc3c1UCc8NlnTwnsdUIM6+fB3j76v
1ZXwF4NmKajxVG/dtzG9O7Cg+9bGO6FbVxB7vBY2PFSfpTqj+NCU/POcgC/bQuD4jjNOfsbx7mY+
v2qJ+QOtXmmmq1SMXzv8ISpKrZefDCYSgMQp/fozeHVbwQn2ZS55GYDWCSQtkbXM2F7nJPzIeXd1
mEGzJQgRximBTSJ5Xj8xeGwHFHKZ8DZSnXphA2fl8OvxC7JWhruePNo34DGZ7dB6xLlB/rAXNIes
XKo3jOWSg+cG2yDfTSFEfra5JoYLc0w/G8d6nRlUuEQHKhz7ZTLNu4nSFMXLM0CNNmXQ/0irp1Vc
oBIP4Fz3OD4mjKByG6eVDLj/iPE/NsSmnJ8FoHvgVi2B8vlsw8IzujzlYafG++uoxyebp/WPMZ65
IiY4v5K9yenObjDAUpnLYIuPWQ8JyZb905WMQmBy5EK7WgkfVp0B7fdD7ETHa8b++vu+9eBGuia2
QCl5OHHLfhCf/CaRCYiXfNh88czdWvkzMfoAmSKWLwWisbXca8ii4v/As+Ay5TX+e58bn1sdkDMZ
y8Pr7nunemLOVfqJfGiT2rr/L9xdA1IWLL4YTTUm8ZdR6Orv9AKbjdkKZD9A1mmhEjfb7+GgWHw2
fWs6+Z71VxWHB1TLLggV8eA3msce+t1QjETvQgrz6iEE9f/9KqHA4JndkW2h82WDxB0Q0xduLqAh
PefzTZZixhvEZEDazPUFvaD7qV71jt8mgsNkHPuyIHKdrd5cOJP8zQgj16SGocC21YdJBEHQSECn
UR/8ku7x7kMsD1KOCnM8Fgo80YQSqeZzE63x/x1dz9N2sW9wa4MQ3DErfOhi9IrkufH3sNA8dkwB
2LCh6Hof2vB4AzGfBIy/2DP8KYpYcg/PiTr+tp/tJif/qarkPVI7J+WoAY/b9/q+LdC19jkOCXG+
fHJNWyGwFW5OYzMhEbqDTBpsbK65QTntGpxHeBV0ceu9m+/3ep5L3gUEdl4NbncNah26tt0shJFg
3agcRpI+Qi37r6dx/Pc6RI21jAS4O0Ny4ou/ZnrjhSyQs1o0Pz+r32vTSLlrqkSjtMKt51or1wTZ
5vHQzZqWr3e/D7BAk6MPUR9k6+yQOa7I2CKXckhCYM6G5klvrN6prkQ9ohufQogBGOVxorxHRycQ
vVUclCykFEzQzmz8osmJl/EUnaRPBXhOiRusTXSiTtGC+zKITkaacEoFYQtnuPI6nXiZSl6HzxmR
y7b4Aus7FQIWrUC28xV8zp2VQd5SSmTeax39SSLHTE4WE5M5iuPBg4bihdFo6F1WeOAbWk9P2okS
Cd+a6SQzDMos0zoWHWpi0KXvKzwhp1QDBWymKdcMEQ1lFb8dA7JISACGNuvff+0ucdRZ9zVcd92B
cg1LxO20XAa5lAcKEuc9Nmn7vpmiK3glJ9+qIxzMCI/EIoio1dVoDEKfg4W1tdBPxYuCsHEyGQ9B
Wz4jLHZTnI0TW51KW+FK/rrJCI5lJ61pfkqQg/WatGJuSX6w0Q3SxdxwIaHC4Gpk4ADs1CNR7tug
0+XhvigXNsAP0Ksmddx74DEIh3YYU6SoE1erCJxqQy9gWnwT0MHTyO93Bs7rTtCRwDUQTWvXkFli
lGDk23etO76XMhkKVwgQXXvKZQgHQYmpabHaP9w0tQi08cdPZKWdkaNjo9sy3xG/eckGhXNWTSG3
9hHD0RgRPn3VZWiiXbm2Ly3280tUm/irvjZtZ22kmdgtQeZHAUW0cTu+kXEkztz1ntE6+MQ+owkO
CkZOibolnm4kClpy7kLYINv8tGsFcI4EL/klZJh9AHuaO/y/ocTnnLF2QcS6K37lMJrr7S4VSL27
9yQ2Gu0gchVVaAXSxTH7+OvhKNxOD9o4W/wUsNLDPNTtyI4SxdClMORuUW3N/3ab6MXBn9ujgtfw
+tIKExXwPv1YvHHgg7MRiAwlZxQkcHwI/bhpxbURr20lZupEdl0JO0EU8KWMcJEjQI+KzQQna8oI
pYAO9HZpORWStTBxYt9GgL+jgny2WOr9ml9YdP8z5xG7nKz2DFLprXnU+A/fpgDYBg+OuTfoOmhP
prSgiUKuqMRX5w/WchatlsJOmRzPEEJu0VfmY+44mAliBSkiQ+PhoHgCgLMjutfatcZ7VATvoaOm
d6gN8pm+nsa8i/uCQqfGOyphQDZKFcpCwIoknrN3vbR4ofBUOC8Aa3odbAB8RbzqFi/26V+vU5wU
4jgbNBZlE0ozdZPxTJRiz3YXyQ17hOP91MjFXW5+QusJ717aP3JjWBsHlJJETIvGR7DN+nmlOoAs
MaAUDNemu5uPoqbXZeBhKrUHct+aMizOkY/Ks0apU/ZOLNwYQkCOjq8lBppuuhQFKjXinTyAVadI
52FHpJogUWiI5Z6gDlil0/fdPMLoA2p4Z7NVuDpAgQTVuaPL/XU156C9zinzmQ1LlAox6Bty79if
AlgC5NEEmx6gfv2mO/r9ogzKHtHmVwG4vGN/AgA/kvIOu+Dd5qhzsJLrB9agyEAIBRN9niMpB+W3
NQJWj9t3e+mlJdiDkVD2xfMKaDIwOJEK3GJogrkT8jfw8IAqZQPfd3C32P9EjTy/lqdEhNOTmHbs
89nHHotMt52ZgJtM6HAL87lhvfkwJ7VQSIBlyVGMZO5ZdHLnloXNZYSjHnVdfR9hawbX4RDVBgP9
ncQiOrTRZG7+Gmex+ypl36N94UIBW4NBmWylEaN3MFbn1KniKijaFaI2GtDDHEV/l+l67GIqzTyN
zcdHOG3vmplDKIIytAkhZO2oMG5RqLkTQwfL5k+2cKw98upEBpqFe+8H3vpcvus+rIF/51YENVWu
xZYyYuaNkSOzq6+WbYTNHxpqeMCF1iTu2hHxiLxCF7yRVNKY7Tz3gKzs2bCttnyy2ZxZCABIYk/e
cbE4rxU5tx5+6bbwrUmzW16yL1RTV6Klz66LhNo0dlDkHSTO6s2X/0n9ueV9U7t9+P5kc00aE90r
x+LdLFJRnyRefsHdPfS5j7MxqHMWhFhX4DmByqkTGSiqrGD3wInlDW4cnP37GEoZCdJHD5A3NAj3
kJCiifPl8ajKBjygqQ3LOAfcoyngPQR11CCdxhoTtSIWJ6PEgFaeu4hdEnibiqQeBjicKwp1rPVh
RbFtBGodEjgIo1xnnvfQO2pSwcGlrEt1Qix0OOTBGiPpyfoKQvcmoadzjMOMaynFuZHeuhHtBTK+
coQUlvlDTiQG9CNvGSnkSn2QeiPhfSj0jerTJvSnfDnnINrGSvVv09KYLeOGG9yYABKuPESqJah1
eiCcPUBqUa7XOhIbJRFEJnCVITFXTQeliTrBFx7u6D7QqzR918PkBARqDdmdJJrAXwSBZdGxj7Sj
FxpZu1NI/z/jCBOHPfBvLuSBZWgEwh9YRuFyJOXwXM8FVdCG7836vVoNKcIEMAuvxE5W3sxH254O
jKSOWIll5E1nlICtaNxO5iuB8O8DXZm/239Ba9g/rfAPRCHVwco8K451d5Iy0FqgEdOgxzp07vZd
/R2CXbV1LHjzvrETIk8/b62d7QzN2ZhpwLcACo957xB1QJ/TJRmAKda+3ln00Vtf3yP0O7ZrRL+/
ELqMeJmMtLVO26mAsUCNCTIBrgv/Qsxdwhmt8cAq3VqGMrxa7StTXJp/FqJtXQQdC2HDKLdiKa51
b7ZuhAWTHAdpynqCzDoDoMcIfKoXzOVaZsK78PBqP/s9CUyJXMiyWLkw9OQInTxROyf4pJy7/JQz
dMZ2ePz3fAbDWWPF3tYiHuKLVfbmO/rkQKsH8jEcP1FZ0cjyPLqoGnEooIN57edVMXP1lgser9s2
Z5douXcBDuaCNYmMLQbV9QeCg4w1nnDhcJ3lbKHzLMB+m8BOjfxi/XtofCiUFSsIofZOL6QYVJrY
KENFCr4UIJgQkybz8Dco0Hnq78tf7a7n6XVmlKZSBkJ1b+K+MdWWvKGZz9BUXiYqtwAuI0Wwbinh
lW+xnMyDrb2IbtZg6BtPvYpUxKXnkVyt3ZHrW9ufoOkNCuWHf2hIMdIwdTe2/ZlZfZxwGv33Xbcs
peh+KuwGSzc9D+9JXaPYPA6kfQIIQRmWndyUSJFCA3BDTVU/kvmWdp3hSKanlp6oHn6K+NaW/dzT
Wli/NTX88TfmeGkBXu6D2RVBL1Npf6XDUm8kLpt4dGb7c8sl9dssJKcmMD1d8ViE0Hchap3k0qLC
paHyXH992LJjHYsKdHP9zDi7D9xKEoI0LSrhrUkFUxd88AUaB+f46JU5frvAEUblks5GcT5czQgw
VzTkgzQFTT5EOQbLtvq+wmFtRYBTvN7n/n4cPSk/9XYDDI28Gn9FYV79hthp/0X38bY6V5Wi1d+h
YtDNjXmVxobzTS2zzuYzfy+fJI/MXaJkGVvziUCFcQt/+SPR8J3Dhq58PiX8dW4KJtopARyWjlMy
7IpinKjR2NDa52Zw+B56ySTO+B4d8cplrOBNhVpbbezTJbFbj8btJIp9Zh8UK65fTgJACh0Iyp9T
Kh7BWxspHtaUk+DsnKXyhndPj5hzSO5fxvUsnzKZBC2NsXI67dKPPBMan+6vKki9GuUREZIVh9Xa
wh+swQrz5lb84/78TuoQg9X7ec9ZmM6rvnHJvyteSRC0wNLS9FSawzUDDbqpn3U8TehN0GcIw0/I
0t9lXDua1Ah46YQHX42l1Z1PQ85Ij83Ek5lfHMHqN2uxZJNWfMTqOTrwbw4Gvf0QqahpvzasBBZL
/uPL+M4jBFqvYiJrCQl/JLCmwzHUPzLEuybJnAR7mShlpjRB1/1EVpk8jZ+1nvA6x/caBDiAIh+b
Acca5/rgG4Ougjl7NRL3rnrLTg1dPIW1AdaDSJ+Ip38oyAB2/FJLz35jG6Dwpn8O0I13ulpW0r+e
P0C0YoOTSXQ1xprzR7B8isccub9dXg0me6eOtCrtk826NwLfe27+gvDUg5p6t5xivtKAZcfoT4Kc
oKDgX2BuB2M6/XrB2+dWwKrfw2rBEJo9Sb+PM8DSHfFEk7auZfQtJkZ8fA3D8Q3PcKcfVI62kkxL
M9nRxmGjgniv90vSDwEcwy2/8PVTjbnAIOwXvjCN3C9chqOBumqx/aGvPCU8fcuO+BHgYY1HN+DA
AwinmQcpy4fVhtVfLeMyY11Y55Y4DTNy5Qq+mA/wDInqsP0YIjtoL028O4mCLzSry98qNi88HClv
uqGwsub5SMECRZQvrAZXFIzvpivk5GdJgp3pNfsZ55bnpmx+TKLOtWt2Xp8qYB2f1CF2U1mfcoh0
Rr6xQXg9ckgrds0c+sG4SsmReNOgdDFrSpGvSrSoeQXJlM+0hlfsu8fFRsrkjHqlIR7aUN7SdwZD
tpJpt761C9d3dqve6Ok7xNMFqWZ2yiotbaKY2RZ3hXaVP1ZtPaoQ2NPiUMkjObyswx9RBZxBSBBt
+SJNZ2jzT5N3j/9ONl1AsPrhRmVSbtI4Xo7Sp8nIEiiPBW2xexq7NuomAKMFKLfCBMBrvPKQ1u/q
YEqQ5cmrMQHxjinjMSq0Q6uyQOlmffq7YhN+ArX3BClb6LcQUYx1ax1kkMNl9Oq8Px4cYtuga78/
id/B1fksPw2LlPXjf7F1EKAHhsQdgrk10MDtDcWvQZNq/gvMbhjYotMDVZqYaC4/kxLSsnkrUYFG
BGc3udCEEC9Mrn271NqwG9Sbs6iiiiktDj/Ih745yFqTCAqY7fkrhNzrjhyvbKsmsHD0gnkn8GM2
ehcbB+5JLgfJtP7h5OaRhkymEwALjgpYQjCpaYTXGcQ+kfm4FKjrkPFy7rNL3A0Ds/VBil9hP8L/
Ntwl2UFeidkMx0oRI71kwPGppPFFBahFEfGBIwwLdD/0MvGAqCBQRFKfnNkUBP84U0mr2XjfMFRi
tFp0rjB77bSDE7Rxrn30X7JThYl7N/nZcsY+qJ/gGyKTgpnxcc4uR/lIxrjq0UwZdMrjc5Gty8jC
rVuRU0GvmMkSktr1V8ag99SONVxCpqNIx5Cn2OvqJne3bMu9ljg0wOnEgqKEjz7g0Fh84AIxCdf1
8RXomS3uw5WyuAWkTDjfxWeg7REtxhKwZOKBTwM+7gdP1YZpSoXD7YaDiRsTQBhcvB0Z03WvnTvl
xiDSSJuzZpUzTvjhO8zWT0apTENJc5mjystZoEQqkjheyJBMh53sWQYA/A4VpUjXCSdDYIG/yZzr
JaLUF8UesRRnF60RE9wyBU0XGAzbtcJxnNFSfpc8BpxvuyDjshbFfucMZIVVqWMsPNL9Kl5bQKtI
in4Q92lznMOkPmUrb/Z/Kx5vQBEEWQOi6ZLaGmN14fTou9eMiaxCqVhs4hT1Yz4A+GG48YuUUOF9
0nfN/DgthPr7/A9LRQlF1Hcmld5aQzyZa7s7WSvfQYQHydBYCpRlv4TQ1HIbKEkAnZYBN8ZrV/e8
iQyUjKI/2uK/M0RDGixsuTkJeZbNKG1BFs7ebSUv6h4N3pKQMuyixp0EJ7KbZ00JgYl92Qf7onoC
ZMgZyOKTi0r3Vm1v59xKEX5RCl22/sMCFoXCt1MkRR81tVpxDwKuQHWeFHtNmkDqBX+ENF2UMJrm
X55EseywF8+BN+F9xNZ71v0SyykZ1wkJS/+KyROw/13Laop4mrz5M5URvkX9SnunSYCBPmft4xd+
qn2gkDDO7FBmVUGhB0yqAZHCwzU8bA8AhueVfUQsRHHY7ApeajaGOFp/nQzmlkI5wxOQPe+hJksl
rIyzRcD/BvwlIRlGyM77Tf54FoKtKRNvprNfEXXrg+pKrqVFQ2TUIDmwI3xymcDEbsCIDaEdIgFb
aSsLi+NWOcXXihmA5jD4ENoxcxQ7imZDghJD263kmqensTKAAbRo6QlSz2L+8vLxOMduUjdxbR6f
mB6s8KgOer12ZiE2/oOsJowON5cRxct/UZMYa7pFfeh1tSuL944NVdNqx3NKuTi5ZWW/eKlgTuo8
0TUGcWHtPZYAqpCbT03ORLYFqv59ohsVvIaYYz9dra3IW/IJgCQLDdYNuB+1VioA2vFwWe3TZKzY
fLohy6i+h8ar622OrKV4uB9RAQzobKwIaMl7gwF4xMWDUgSH8eAaXzcsi+fxUS8tkc74wDWKf5/f
JhF3gZIgzTIGNMIe47qIYao4zkhpzdCdrxJhGXm14L5tvQFJUYtzvtpWNVcEfLkognYXY3Nmag9R
MkCMEqujPX0o3jPH80KQiQA3N2ft4kLPWRuTc2LpHPzwxn1XOzjNhsKYC3y3tFD8CIPBM5Co8HLa
5N4CtJEiFaYXXUANKlOmFHiejvdpR5DR3Tpg/LZvHmc+d4GS3RmwAYi4+2d3+bNNLKLpDwHLFpcd
1wFRaS6oncToHiOf5+aYWxy0dT/iIzAhedrtr5gDxMhgkaY/7UHgoCKm/tH5LUMHDL3+GiPQEMLD
ytC0hO0Buhz4dHNZg9o2xdjl1ur/Y27MixEWb/eDWHd1iRgYf2TKO7c2zTP6QBjqQMH+7jr3pVY5
JAQqm/AgQKbnTYXXgrpTIAL5/eNck3HD7eektqiXWdQWWD8PCB0zQJiEElaPRAiex64mQU6WDbUh
RDaC/tA15iTe1Ao0J/wPleeXORyQzA2nrJ7hEui0Ov5Zybd5JAerZoot+Gw+cQ9rXtDosG5PZFAY
QaCm4IINRtWdfmokpYQIIICwe/laQaypgSxFCNg6cAF3FNfMACkmvkZGAjCuxl/WMtRBtggIEj/R
doQrhheGkNXUYIj4Rj07fxyWmZO2mO9Z7ANji2cKRMwyWpSkN/OEF9098uyNHDKaWYG0nj5+PyV8
J7+QB+cYLjofMtFW5VfTJILJiBWPj0dmKvXqQoIW/Kw8H2RfovbTk+SU0QQAwAewmUEh8G3dHc/f
DBEczz3xZ3YTf5f1xGJ3fB1Tg+NGjyu2+ZDLK3Oe/jmqd9J+7SbHIxOPMJVRz1hykj+pFxMpwZjw
EKsinDtvVcJbDbiRNO/yHhYG7kn6GMu3P3SBIcbQuP9u9LEiP0omrMVRBt83b9xW0B8fipoqTavN
bR+jw7zd9geQOYflqkdauq3/sKZ/37rl/aJnbuVXpauBCsJ+kAFfdpxF+tc+yiLgiNHziNET6Ax6
lTnA3wbNSJQGqSBj2n3pyE+1rSeQRD7KE1gK7Gtmzn6eonWvwAmqzhQM4aWS/0TnBaulRHPcVz4b
u50RgwdRPGAzD82z1UJYFymjA5gZ4OCd0zZEQU3hPEF1uIc8n5L+jWwX02V8j8jg+1PWda+Lp4ug
hHop+/k/zvR38kF7EV/IMoIPnsZcq8FwA9bSAaudTkem0KiC1tz+cpT9DkvLN3HtZwduguNpdrR5
onctNx+A7Kgd+PfR15lSvTzgM1rJ81ZxU1C+8sKVePi6axB41a3pyWAqSIp5YEiea0rmKhizF+ni
ljXFFsIxLalMIxUArhL0iC8zoD46MCNAf/wRbbNFXWL71ByRieHdsJ4l/NxhPlNBXG8Fx7Alqqp6
2T7N23ucCnGrUq+/YXffijDjteuRLIyGQe8vspu8VLm/14DBDKpOY0I5YEuPnDPsYljBosg5e9qs
GZN4HLsxmmsdFKznXyTO0IJbuSkKnasD/msXf3YbDmOQ6z+3niHA3dsHZpeFkqWvFU9cQnARtdHN
vK/gs6WijxMfckibXRp4o2yC7yL8AAsqX4PE2ouNxlnsmJC9P1Zlkf3LuJ3RUIn66mYBWfWHTW0V
miDXFedPisKScYuWIg7XnHNc/+K0SGdFi1+B6W7pmuSTH9k320cy7RF4/ZriLBALjDj/7mmSNNsg
SKL+uapcZfP6wWxWxwFWEmOdWDoD2fGsOUHNLrrmogFS1KNJ8uuxwxgqp5IR41FJ3puqpNoxo58f
1pEzp3j+WX9GxdORLjVLtPBtOa2abGBTL41qOuI955uvobR7V3Sg637KbGHJKTX1651wPNhnAlHR
/d57HniqmGAxMQWtHEp9x+KI+mjo/b9wYL37q49vU1EBXUf20v2GVOhf+5nuBhweZ8bUtV8WDCna
rMf3Y9t8p8RHmfwk8tuQnkLH/QE3agdexicnr7J/2N5sandnDdytqwtTJOnUCZ2/l9z8L18XnhY6
/NJ/mvlMqNWe8bAO1knJ+AoZzvVo+NB0i3ORWV1T7uVo7hnsjT13YWlumkWSPhGLc4lmLOiBt1/K
biUbC60wSZIp+WNDFXOy4Hzw+m8rE49n6W1BCJLyCF/9fS9mxUp/BN5ySb4bHL4YiTVKBYXPU+ja
R3H2MuNqdXmL+B0VOUsue10BJMFxc/Eulr9smhxHZ5hhToKRuL5lFcGQI4y8FvM1ewse9+cKFVmf
WY+H1f02LMKBUcmo36OucjcsCFNvQXKnau9kXk8BpeXlm/A8N84bcq8bQkEC4pBCZqv3iWWj0xDg
tAHLSXmjPT67Y5mpE+wf9euDg5bUq9zjpbpbIStuHpBjc3k3Byk3OhAVg+vIjC0MaSMmWiO1pWX9
gUMnHOR4ArwSzFysWtnz3g3gK2VRMPPIu+OyJbLwwETDidb9Q9kHCIp4i1WbEvqo0EpFS3OYFdFg
oRIPiYeiZXBwg4FPpSTkwqeQOpIpBQASIIoLAMX4EV0e78L3SJDp+YGkI1L+Byt0zWBzsjMKUa9b
fHYxqJ2uTcuD71zfii0zjuhMTtYyfm+guX6yLNl2ZgjHIy0Q5zi6A8gvzz6QGxa0tr5nTFh1IKg1
Dctdsr9EJetKnmys9DvhrCx/yx18r0zKR8KETqi8f/+7UOJ+xq2MDE4k4AU/P4imRbyLIdzMZE34
kv0ycuayQTDlAtokaLD+VI2GmHvwniu7ERAN47m9S83gDmoC3KQOBoP1Ym3bosOJshrDpWdCAeC8
KFpu14BEWaJPk9RfBFEK0Y2kCHphPP8G9iGU0yjUnnEm88aVZrb/bd/+EXZQWG0DG4WAxCq/R8Zq
4svwMscJuYM+P7zrCnUil3nIstUVxsgkKjRcOmg3/qoixz+0g8uhb9Rh1gWA6yJKaX82Gb54pHsO
mVeKEbwT+xfkaa9rSzDinXrVfmwSmibG8w1RkYExZ6Dh3Gqk+WGWG8W5Qpls/82tERYTQqh6mUM/
j7TztwUlY+QqBbTjczuEl6RZFNC7aFuouf0o4nXvOIcWU414did/tbxYF3N8UmO52DLp2Bz45iaV
RESS+DLQsUuLUb7ofAIklPAJMEYesCQBU+Zrsmqo4h6i2cMtiq3VgKzL5zQEzCEdMWuFY64FkIUs
ZOGHUBNPm1D3VN76nccHgIB+DvLU81p64SZ70r3SXkNhOQZ9eaKwC15CL+vEZvXXqPc6eUPADGNT
YLM9xULUkWarvSAPgO5fzwkF8O+TTA/FqE+iy9k0E1WPKeOxRNMQPCjy7IM5qfP1iw3EM48O1cs2
TPt7Y1JpG+XXdN92HmPxgKsyWtR4fZONrXUKCFTteuOwB+hYp/HqPAu0VmfDoHMLq4ebaJPQ7yAX
mb8a8Ts00zWv2dSKjoHOm97i8ll/AIF4j4JvtyW1V7MEByPK/n4cHzT+qfR7U8KlklxcICqjESxC
dw2NEsOZDi0KXhaFkAWy8kwbHD7Cnb+ezrKeTf8oDI1r7ZmhNYpRtfMj4gVFtRewZAkTq55giltf
CUqlZI6euUTXSs7wtzL0l+plFdZ50kvalMb6ZLfZYKLh+mF6g6hamcKh0H02+WaT58EWVqw7lgSu
J6nF0uuK7D3wUOA2K0FxOmuS8OauvHptF5e5CVeOwTSkfLp4W+Ysnw450dl6qzlMbh9P0FDttcWG
fqPR8MCcAkxs2m4/3Igv/UpW7pv696vsEPz3Tn2ohsxqMIErIZ9FSPNPTOrEJSjYKmX9PFNyw7Kx
PNsj4NFf386dj/YKmcJvIr7FGUDU9AlYIne73NPg9Bs0r7XMml2iOedoyi6BqWykiBbRe1N37n/9
iOYYHvF6hTAg17ROSQV4rmd2BulhVQAxfY8/NxE7a8LcYwoztIKey0PNVHZ7N7KfX58qx7qYMFCV
p+7D+EJHE8gnWJ2WaGSWTjNfsTZ/a2kPwhuRh9IKRMDPkKXhySooOjvhFaC0uDnoz6TMrWUnO47I
wh32Ni1Bg2iTFPZ5bu0MTqMYNanpR/7ho++tcB9oe57s9shdspYwGAxg7W/DTR1e51t2bjhySp3N
MDPbAO/plpByjSO9RMcIAFUqA4NRTvNBgZznnUoTOblRpE2mvH27THPs9F7KKnxZ5xxbTnC7Sl/u
6Qe4DgEqOXhDKJFaX/zDlITOa51EjL7FbS0z/M9YhfgTPNdPVg1hNSGirrvNX+Zdg+vtV4lkhfjD
Zw2WMNPl2cMDQegJM7Ku+aqqosBCB4yAWNIXZ6rWvneVTYSsbcc892LrxZXXxKSmRO7fImXH8MpA
S3kWYoMihd9KEbVoLEVzv1XKOp6mmeWrSZzJpOLBMBYV8vU0XuMu3ja+yRfU5SFKBIkRZsrWJMt4
uKikgPGDiVI1CGGWg+E48Ue0rwX5kV0NhYXFX04hzHUI4lVLvzc4ohhNe8meqn4Fu+d5vwodTqfl
wTePCQylaVIYRCMP4Dqz98sb1mMo6HThhU48RB3B2KfgYTyuud1ivxwwoqj7QLNUPS9ttHdBz40S
ME+9YEuhATecesh55cOhiuiI93YSykQWxAR3zDlwCxpEG6Rn9mMg1RZ0UjfiCHnTIHxMI8obYTsk
culowTSetK7/FCmoUxG+MG6+2X99aHAI6D/Inpaf2BQN//xBrXHLeX/vdfg7t4sUVsw2oX16UK7T
fJBsCGQMilEpbZ/ahAYcvdl81Q8QQME5eBBkmyl5z02bu1MBE/eRRCmmdwdIXBP+C+ZKVludqr5F
Rbj6BJIEKK8SfLSoUyqC2Ws3HQEIp2OpufxvBN+APH//U7GSPSsK279nHp9xJAPWmUFKFUkiAddM
eI0XA9Pm+RNSHFcCx0nfExS6i4UTAygpnO9NMoYXRCs5YxZsctZ25q482cAEll3GK9uw11ml1AjZ
Q2rKZJf0rhShLHB5rB4LmEolKM0CRsnpEtO3izFU+Q+nVionbuB+Xw+g+0ZQtCykRLqn4u3h3FLf
Ct7+lgmFvtUHQJxR7tGXzPZISikY8Z2kk8uIBrKlvgl12Pdvl+L1QK5cnGBa9AyGCHSsDCNSXI+a
N+o2gdWRaXQwHTT4m1gfts57VAOCiwL07TzJQEqRx24ulJaXwlvzqIz8sHfCWS/xN4T4bTBRX7Hp
+28a5lMXWZ3o1clJjPtGVVYbyJJjqZNbRcRkeX7LPux2gcSw0BnGE7CR4BTsox83HnFEeTkYCluI
HdSdg4Y93Je68BF4quljP/PS9Wr+8iIyiGcGtsFUCU+Ct0YXZGXHIFW42ZawKdV01R+03gTUCjq/
7pQilTK3bBpCJ6vEQcujzQypEfw7KzpuEI6jhUk5MGsNmgTbuABt7gu3BiQ901gPyPMQd6IOkjkU
rWAEbi9OkSWsuxfmuzBvpJ0KPmc8Q+yAyndIuu7fNcoud2KWYXSZMLeQxtdcxKF7Tef/yoIhztz9
lvIl+TAKq2sBDUgx0xanGmICUGphhNo2+EWqj3La2mk4ERrRj0J9S0LogK0pe/Cn/4+Np2AUitym
xx/NTtV9hfxXwrrJrG17yq08Ebu5KzKGX8kGrbLgftU6P7HBxNQIxqP97VsG6Jh/XbJ38c323B/E
LiNHIz4Rawk8mzCVuhC2wtyXjzwCBfylSZS+Ga5cAzo6KrBOQpJUlcQLhsQWaESuu364gQKLHgtL
acJ9m2qiBZ5ooArTJGndrtyCeR0n2UzeWO8+omTcnegLuHIhhmx7wU74cCUybPUjABP2pyOCQ0mT
jNQw3mjgndEVXlqb+qsgxhkPF7u5XlSJxkA9a1hp6zXOEf48QYxqidABT6+ZERM6BzdhZDawVJB7
yXq7E4lOLIodRq6mj5jCQZrNcodad4+eNGO12zwPGwy7LEIbV3DDXq+UsEVv02h3rSMi6hBq1NTo
+hzdKttBIhV6teX0UnYKtkjUDd70GQgFxqsHOgSU2X8zBc4i08YXU4ONDhPkmEpQX1q33cnVxASL
XiNnWb34NEwf9hfk5FR6tTKmwm2n3qMfsobaMjYEYKZ09QwZKU+c7V71XBQ3Dw4m6jnN3RAzRIpR
5aqUk8A/7bBXDOkGtlto+8RKzB7W5CisqnfqiCVHxRnAJZTK/1MSz/XafPjUheZSXnPnTMZcuS1L
+nRCUh3vNAoZwBmdYN+D95eAkVERgO+qLNkbErnjf2OqBxpv8vOTq/gTtOLtZCqqAIeT04jDlpUu
5OqV82RAfEZKdmb+QPn0gJx88jqpoNu99krQhqO8X6nUi27aJeUHqmMoI+Hc4ZcJhu7N8I3c6rmg
3qvcO15N25POcqET3SosmSmX9LPCj+VN5ps8GmDsCpVqqMKxQDmd+uuSan/8LkYlDIe55auDg3v5
wVNVfd+5BvNRK+BeFJBcEUGMzqJNFSc7FhXbhYQvMoOsEosp4WDZqLmcvU2kMoGZRTqqFmhEKLjO
DQEuJ3mgHRTMAEJ1xAe1dITMU6LYKystG0VuAXAEugAgI+f6QKPc7ijMrxepOP6b6OV2owvxIsJi
bAj10CNqG8hwuPqtEnorJQPdHhQ+0R3dKsPBa8YsTec0r11NU5scg5mV9Cs8HTVTkSCRTxW0/tI+
0AIWz/zTiF8YbaqG6ipqnvtLCXBpGdHtgB7sim8cmHmGYbmtOjKYKqw2KdppUDNlX7GtS42DXPJR
wPZu+U7tB2TNRwMholVXNpm77X446sdNHZ49Y4zz48WygB1OIw/HjwAqysGUETLzF7a6eOOWYKoK
XYhKw/KyckD3rb8kNf9d0LEgYjCYZSicOwHT/lH+BvMx4scYbI1T3O22GhXuh/cO3b/cs2JznWdD
RovjHSXH94EjRlmRLLbGoo2gohmzJj2Nwe4Ktx6eoZRHhAIoi50BeaRpTGDteQSk+quQwXvu/JQm
Bv0zQWti4M1S99yRnQ56RDKUUMnDuJhbFniiRlIRxLicHiO9mo6+rPRu6mrXzwPHqSy2gEdWWrtW
F9roesDmzaIVM5XxyDMM6EhjvzRGlQuzpkHdzmx50YNHgxwcHtQhTO/Y4g/8qauJXaFoi/HORXAv
rYAsIoEhlSpGbIfV5SK1EM7dzr8AUEG+1UhZc933UsbIXynMyo4FsT1RsQOkg8kDNdUXDyqzQyM6
+luWA8D1Cug/fu+aNq4yrsSCOw8WqMJpP53OVpx0l2SA0hCnQWPJDZdTvFzWxbxsZ5rif/HbX51P
M4RlGOqeqn3AKnyetL7NJXZtqQ/gtdO7FzQC9W2v3PZRb8726rL7fzkrYcBvQQs79OydoPfnN80F
TvyuRaY4DI4i039SFOfpSg6MMdaypuZh9iEyWaOJniUXuOe8GqSMmkNn241Di+5JtAOlyfkY45wy
8c19uBsGDF/9jLNuq4aoWIVn+zu9RKp0tBiittjWCQtaRuvfUOyRWe4ZegNCWBrPevpm/NYu/M38
sZl4O0um0hoNa48gyJCFatsYOU9OpBy5Z5jypWWUG0sTXBg26qaMnSbtr0Nla8VsQ/qSH3vZF4rN
gc8c6buhbtEA6nJ9XNF7DwaCOVUYfromdvntBO3WJfo+1IvG4Y93tXgcK9ZSZXYgFbzHHY3gNf0r
9Jx6Qh9le6NTnedo2DZ7JJa7SCKuDrrJY05rUvW41xWwKSwhY6FZ+jhcaOMdY3L51JpdGVT90mZC
mfYAi+XmOxTwDutYLaLJQN1FbcALFMy+oEtXZ+CcPsNWzmAB22W8BLxsJksr9///i1OjHdox2GvT
VYgt18DXSHHUUYHKCMBdGFU7bDKMhn5ffEtwPtKVzpOk2q8HsfdcBCbz9jV2olplzMhM1akideSt
/EOHIWzycwsTvMJDNrDxSrVzU93UdEg3xXAi1gzoWI1vwsyuiTIUpfjKJ+nSiFZkHZ8mMH01ucgP
3bchOSDvJlcRqlFDgnu2zd0dHjkRR+CZVS9NzAbzi+tFHVxyIVesdNUOFKluqMa7D50eANcoLPkI
lF0b11gPjlurbnW/hzWOwdKkTGypVRJmhXVk/qtyIgingm64QV39dtVjP+1nysuZjJMPUjWd1KKo
oDKQaA1fiDYJ7IaMANRZs2K5xmjAii2M5qxvmI2sRbEj0tjYGKMEKWuK80Fl7Di8fU+N+AZLB1dJ
GYTsH2EWMQ18SUdTPVZxP/JMS/UNcaUeKhs3HspFqt5I99Irk9SbVDcUGVG4gIjes79kApdZs9Sw
fc7iriczxLxL7RC9dvN7dtReJzJ1AVNi/CuKZbrxF2q5NRoAnhRQnIJ7BRbiBmF22d1amQbK0aCh
mKQiVK302hZ3Em0YnPI0opMjtnXGx8KrnFyO7JIZmxHFv8Fr6oMNw6lUtnihVAA86odzrdi/scgK
zOd9bKQ0m/KMl/FFtd9f0tVkkxrKR5R3F0+OSpbfvJ8GGR9K4lNRuO53p2dHb384mRZYr+goqGN1
6CeuzLBTyJUeI+dmJd0NHWL/35kISwh740NptntMmRIyBZEuKTaoSpoc1LINrDeF17fsrNkQN6dL
B8Z73P+P9iToSIqNhHOMNx1Z8RkMkdXsbj6AgGgZUYFFciQ7lJiFswc91jjiDc49kR3EEdrrv0/w
iG4kHUFjFxWzaTV100dBpNTv7Kgj3HOXOERQ3iOpbINBtfkv+Tx4L4WP39kL9zMKdcorzgD+DuLp
EghB407VnA1TR8u2m9iAurENlgxNSWxN2xN6+MrAo3sncz5S23RS7plVFkkHIY+WX32bs+ZbjHeb
2PXl1qYjSExO9Mw6Q+5x47LFVvhLTB0ZVXEKVB+jdYxM6ytXXYu++pRUpAb7X60EG+b8Mgypg9yc
7tUkSUP9v7H0YfXxr2G9eHdd1B7YRckRHIUu0dDZ7NGAmD9ldFUpWI5bf3POaOgEkQTpdUNpYeUW
Dzqpb9PHs/bOdG7b9c1Ti0sQTSag8AoDrGLXcSs/WPIHB5ADO30Ndo/7snyhq9L0FEbcGM3yc+sm
Sx1NNaMD4Fywn0167tq86qjTxVHOX209cxzgp3rjqk1nEJ1jl/PosodhX3KqgovqE2ONfbJQ15JA
J7RFyC1o7pFrQ+dSeHe7xi1MRjyMC6CFEnhiUr/+f7dlPm28bBhaKupFpoS0vNHeSNMeOR5PslCX
hbMfRMdUg1d8cjOELasUiPoxP7A8RfsDheMVGKKui2H+t8UieGgrEf0sE3S6Q691IuyazwbYIMr4
y4scsiZfy/0wNPYXAvMY0Ge02E77WGYTat6li0sLnp6SQ8CcIyO4+WS4tufgQPTg80fFCDPDx9zL
D/rcA3fP/vZK2gWtiEOjE8CPquKgOLjnjqnjr0w2KAu3IJ7vpsmgp+V5aJNeADVXtlGIBfsys4Og
+AKDIZzwZhIgtsmHkcocHZQ+06UtN87tVx3cKNeHeejgGhlI+6YSdQZ3UiNFtquNQgNZSsStMUB3
ye2MpO4Q3Gzdb2dvN5YtYZjCAu9JjpaCbgOqEToF8NyY5k7SbA5GdP/NiwYMMgo4DUUqyH3/D8bJ
pamaTrsonFEdQgihk7+uM/qGzTYbRwMNgUtQRcJ7ugvS7dlPOqDVhhyd1JcWwzUe0DRAakgvHMGr
YqaB8e33Kn1S/PSJGjm5GZpSmD3xC6vI2RNcYF5jaztvuSmOlRgcGV7gALk/DTTD4K/0ZatpRKiD
MVxyG/5FfDavMRlATd0MyRXrEOgRxJzCsXtIvYTtK37PBLucjhr6JtFL1pjfYN8daXmRoosm8Lyj
6gPHGfHk2/uCRN2B3CihTkI60kaUivjOpF/YWxGLyIiVc8L2IvXVjjypxVBUmo1XOwRVlhcSUZQC
mCmNCYgyn8YXk45Pv+eZXv8WKGiW15rEp14oouGAykp13M+1ff483tqRDf/EguHXWUdLpoXBZM0E
fkU1hZe/NUv2DOTiQ0f8gcwx/GhwfCkwZlRLChGf3mj+EW6sT/vZx06Gd5PFqHYMn9FrJ98auuMS
3TxG7LWTpTg4WqqtF2MkWabo1eG9DAFm4IjEUEIA18syGnl1zYzju4KD8/fkIbSHzh1Ng2TH1W6v
i3dmWEaHSlfrk90oJT2+1QHNPDPPwACGORH3Jjwtfi/9eEBFElM15QuGFwoKdN4Usv4unPxtyiIr
ZjCa4MHk2n2AenLXzNoiwsn5IDPFkt9WuddA6iGlfK4kae3+cPKbQtvtDxrQJqDrbfU/6NcT2jU8
ClizfRUrHO/G+DvXzwlmqZB/h2UXwrckyEdMU0ty7ZSy0rcLS3XXs+ag9iwf0Xgs2zHC9fDJ2v9i
dKONCThsdFNhPAC/wXtej1P8fad4sL/ublGhN8wY3QE9M/qLlob2LuVOPbXVThOWPDATrQGWi1OE
Dr17EMLCUrOhqb9ZiZ0z1QhPVBlGp/yZq4MlYp7pGv8hqzv7IllflLmu36i230ixBprH476AvBsJ
K7shqHwGM+fJeWfj/Z246/HEUKgP2YoyKmbJug98iFzt5OPygmjPQWoE+ycTrkxJQlSmL6VJy0aG
swogjtFvU+Hqc36oDOU7OW1oZpf8xdgEJVNBq4Cyujr50Q5M0qjgcdrH5W5I0xPHSB7T3E27Zq1p
onuaz6dzwsdq0tYqxaXisg1BoE++V+QBAn8uK82gJi4nVWWZ/xxi72whYW19nBeDWA6l89DGb9Ti
w4uIETV5LJfnJdh1dA+WuqZT4O/khsU2rO58GLAfuviGU2j1ZuuP9vVOuWVAJpV+qEzgl2jVM8x9
yRgP2139WQwJ9wiSam+k14vWIlvPCTnGE/a2cGGy6uKDSYRANUjVudgtI8EEM3bDJ/C//jTGcWV4
vwsytAWDIr6r2hfwY4ZI2mW7nNubIojuJabllv7oRnYWa8vV8c6hB+KClOCoinh813iyWTX1yXEd
6t0Pxo78fw+yC+bdzTtSu4ncb081Gl7DQBrlDo6nmPpmuEdlj7ZkU33K+DxxDpm8S6En3sJkNOC/
+FOiTlom20kA0tl6FNWylHnMvfOSeuDDc1jUlnysIoF0705qQvKxFqybjHMk0M085/WI4LY8rxJc
5zhRSvOYE8kzLBcHJwHjpwa+5Vzr/pN6nA4+Y7567laarc+PYTfokXt+aifJalYFGpVspoa6+ENV
YIqZMZzqYPrkxH95DGNxD8bITCznJsWJcsFFVmmCYLnuOe4jhe8SUNQ9ybbPXg5uXroCVvsxJ74R
HGgIUtv+WkZf8+xL/2wJxQ4n6Q8lccTHCl1SFBnE7xIrXG4oJOWxnWg8cCQNz40Le4tKAzFF09P7
o3STTEU+02SPYx3QH2IMO96LdnI6yLOy3I5wxaGtDTzDHrsx1aR6qDSumWWRyEdXh9Oe25AKxUo4
tV7sxWkfIjuR2auFvVssOA7dd7/4KqSy0BU1bEQQzunZUS8ETIEMM4OK7sXFyc/1gnzMHv8LkCR+
K6jzr3jJ/4F4zYYC2ThwcNV5xojEdfnPqlDgT7RhGrwyoKhkx+sPc7m2UtIAV2OiIDlFBd4bCK/f
RrgeD+kOpkz8iQZgkVJsMrQiQWPcQKuUcK0UX9kPseMXsAMZ9eYTHwwovfPoo8wN9/JXR831NK4a
cGFqb4dvq1kN/T7U2NzfcCyrQsVacHC/j/GxXgIN9AwkIPWeyYpm207dQ09o/vYPkhTCB40uLNXZ
4FWi+UrJ/e2AoBNH2zqX7mbgmrCqkgEyFqQcYehluX7Cf8C3q4wrPUZ6Mt2W50gdGz+lCztMdt0v
FFmtUUxm6E/atlMbuzoSOtTi+wwmoftD3psXAPGviZs/eyg3QLc0JTSjBlfjM8Kr2xlbP1MEh0B6
E8CUUUyChd5kYFPtjMLvETheR5dMwA70uhVcsHficDUSG8+Y4Y8IDk5X0tcnJLyWJPQ4hIXKroT3
5+LnnCtYCWD3MM57M7ed8xSPJ4BMp+UkA3Lyc0SVItsb4OhIquHJUgv1u2HZiwE8IRDyQJe2YulJ
V/Ewe9vp4UzM/GvdLiK0jz9OJgP4WjGcFv4LWcgYKqAIYi5mtDllx77iCUTMyxi3RcUZLPQm+0Xi
aGOelZ6fLcbCnNFqFmpRPewl60arLeVGS8lgm5FkXmRHg8Rhc0GZK5rtacqNlScUZlBtNfR90aQX
Fm0Pk7J+ay6HaiWmWSHAGUKGnNMwJo9LmP7OAygxI0jhi85zPnHBO32YnRT0PLQdGwOLUaHp9bqf
7BBUZe8q0MiYPRGge08WWpNt6WlIgcOCRoYdTf0qiQ081xGUgQ9+tSmjvNWPnPu1xuEQjtaR9pqa
WwPTGp6NGX37zdrJnMqnwAKQI+L6L925A4aV3zoPuF7ExRT75fwn+85Rh9h49kU0ncJbkFOiB86h
iF2ubkiT6/rDdT5hYX9+hr1H6P/5CjO6+WyJKS02E00G15zAaNGrZA3cMuMBM6D0L+nOL1VHjOFG
jHwucxsqLGFkZRK9B3AiT/p+3X/2DfCdzFqfly/gwTnsxXyS2TaK50Sf1V8Yhwd+BIQ66vFEYy2s
bNL6z5W5xkROuNAXzNzCinan8BNxNnvEOHMtdDLo/rHexhCMvpEGMELpwhcv7oKmQ6eSAoKV3Ppw
EZ27Q0mEMdsHX8Hi2SgnSwlu4VTUu1cJfRCYNjQASNMXl3hnju9s/9ENq47+h6t5SZpagcNJGV6B
MXmz/nEJoDziW2kPr+KE9xd1f0w1/XVMWLKqbsQL+y+X3zTHi4UsPWyozB2wSulJXE7eqTdxUEnE
MVxjEUMqssMnx6Esd1xxCWhfvtj0jKqXMwqewkPA8fsX0f8r88ORNnTvmtN/Uc406EEg4RGUJI7A
JjG2eVpd96EL3Hkv3gMTXglXnepx0VML85W76w8pjPaOk1/xjXmO7C/dOKd4eZu8Err5hNaPznid
bZhh/StwFNGXN/f24me4jB/LXpKjf/FbHxId83qGtQec3dQdhSY5Rk2YQMgbEhY7ceA3VNjrRtLf
sEK3VEdKgtnpeb6rrk9Ab8kAcEjfWK7AXwuAHsqDKKm598FLaBMD2hGHs7iQIjseCsnfCaCOkWba
0MKYzeDHpHWXuHBkDXlQPaMZ8uX3I/ixxT2f8pnmRH/jvYFBrqLuSyW7ejwHkIsUPGJ1TCLVxRIh
CPUfDCX53NFmiWLICkzI2Jx3FokoiUl8tmX7rKql16bwTuSeqwYTQCgHJ+3q+QFDyZibfyi2i9c3
NpPDWdAUBseblhd0StHG5pOA/xAALW4rP/k/dUCCLscBmaxitJFegMeKvWwv5sv4O7ROTc2d0p1m
Ia+WBhY=
`protect end_protected
