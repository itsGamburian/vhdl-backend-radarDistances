`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FqsgIzh+a+kgdV+2K8GPG0haHBTWy1nYhlXFDgkwRRc8HFVg17MuCVhFO7CdVF0qtKi2WNw/dXyG
2vqzeNo2Kg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CNXxkcm5DL4NlxBtfz9iR14F8tJyLabWEflzi/TN2Fl8DtI4CFbxUwUrh5b3HU80kO3QFwI7sD1a
PRmuiZdlwXCKnYp/HfVAntrf/pPawlqiBTXh4/ej5/bI5CtdYXfVYTa7yPQm10tMAUt59unxqXZZ
QDTgU4PID626v9Mqbj0=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1XBrWt0OKzKUoAM7/1MlzHW7zwfeh5crGE/BQNrJbDk35j+JTxzp/vMXc1C4AcpqiAWRoMYieUhJ
qO102rgl9PNIBOUva7mGwwFTeNw0c4RyyFIOBlpvrRtnL7wiSe1LDGLiCbyQgFafxoI7/FrPuDHB
h7eWDt0u6gSy7wIY4WU=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KyTRBh/jQyl0UNwJg8czZOue32n6tniMI1D56tpVCIGRMdDiiOrxhQaRxp5cQPvTQ5PkOsXqaBVl
g/ZcSlX45jieea+Sn3gIEuwSWbTnRwx+BLyCe7EG96HRQEI1UugacjzB/fnWkBNTFKrv3hOFF3hA
qlDYxrOzEboQGZabNBhcepbw/PchdzJThs+TZlNR2aXJAindqnMbIC8/PuxDh747kZGPlbt5Pch2
7zudV5x7yQlzNMai4EqBfOvkg0N2u5PEOFS5mVHaPVDusuwrxy3DQ36fyQdWhnsKaXP6Z0uxowV1
UROhQiaFL0ZmWxOucOuikCjBWMKaGoUEzppdDQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gw7YomMKO9TuPvP5KVEp7DF4CLPn5IjsqsfPl8yIY8cj6JNxM2oQFamWiylh9veU4eWC39LXD905
eqMsuK5q+Wk/FTZwYdNVbPzkvmdSFUqlkDNrzVP9g1N4rnndiy/sBElJ0JJ8PbekfXyHfH61oyj3
yECZCIt6IU31EaqDushYuB13mIDKIFf+15IQV2o5Op0rqUXzUmNh5JwWPLvC6xRmcSxmTHGJj44f
+CbGds+Y6NqiFWTSawVmACdBzd7d88fqUZSUTGp6PUGGyLEjxb5JzzVw4R973C+hJrKuyy63MtMN
FBRIDs3/QNbA/J77igTnwvJ3JrINk3I29RjMkQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Pgx6c0SyERgsEf6fblVyjdTWj0eGk4nvRl3wQfTvfIZN59DFF20WlYqBXLnDawz052Jhz6IjeVRY
Co5oshyXJ7NtNVkda2b13uvYqZKhRRC0Pp/gdz1M/QcAO6nnnI4KV1ifa5gypMsZKNxAZo87/hfh
lLPjL0vwRHWvpgljWrF/VXrrP7ZJXyNXjGJ9wUsk7AlNNUlezvxMcsoUyMgraY7Q3CJPWUrgHOCm
8NCnImGLP2IZKAuIcC/RyAkyckR9iyOX7UwM7lhuISyHmXExliZxnubh9g7zARdWNQpEoxp70a20
wwDC03NwA1Uz77TkahUublN3WyVLjgBpUTDXjg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 565792)
`protect data_block
LyW3vxxIXyAQ7rWhi8WdX4hJLWCZG0gMCPztrkOqpvL4Dt/SqGz5y3/ne1vKOfcX+Y8FVVY7mXys
rnR+JxMbwA2PV2/GsADrBQEeSdHHs5Rm0+8eilUTgoJdy1rj7WWpZhGo95xPS0Jl1G2Hm9crDO5L
bfRrzOlhCu39TAFAl/mHGviNCgqmnS1PlIE/2M4NGlXqN5glABfKBJjBgXyMlD+69kuUfvzzWG9l
5GgHS2XrQhI3fRykyCUSNFLCPrSWznS16iqDihWLaAXc4yc6SWO3wvoUThWJmR0hNvop8Pd5/J0k
MZQrlmID22daKrgZ3eg9H4Zsnhsz9/pHImKlEljEKPLT8eV3GkjG58B5O6e6OUtMli049h+OFIyg
/Va0/Cp2+JR+TnJ4l5qzAR35swSGAaTufC4jKym41C5zKZNWrm9B8Yx2/nUr6HK83xmLKNZ1M7jZ
3zQEfVLJiaCyiBaeaer/CXNL3QQNybVUBgGKeHpXQAnaJxD1KY/a4EPvMslqQuNQb3AuDSw8kJqF
e5hAv6aMH+muDe8M3XOeXhxfB3RxlCe50JGtPPQC4fCT3f1+Iup3xK7NnvmFKNBAy4aTmJQEyYJj
LFwToCQcFDgSXdkxsTrYm45YA/gun8Z84QL9xA2dTB7bCh1JjjDCqml6iTNhEP3hLFRBRLHpeAcp
2++t4CKm1L1vbJykulA/oJmly2K6HMTne9ADdK0Ytj2si7CFQSG3Y5WLS3jYiPQF6fo5NCWw3qeD
Xl483VqHsvxrYk687q8TPuX4enYj1Y69PK0tsjcDCtnCCnQiK7H5E928EmI0XDUC6Q07ng1dKMD9
ZumQFC3UsFf6AUQxv0GGntfVQ9/61T8s/kEajzT4CzRRME6Lxd/s2rPVsHGM5RT5v+OvAEwLz6bT
gno31xtusIVP+RPu8IP7oaLGPUUTS2MGF9CuibKDk37YBOPPXdv93xKxr8T8DyqsAeEFFYT669w2
UTHahSh1evfnOGQ3EWjM32YJaHFNsjiJBea5RKBJscYAakIMOKDz5oJxHiPj+Ac4iCUc2E6rBcUU
TnTyiup49mwgO0JpTOlPXYkobaj+2GN6AhMVzSJ32A3Jxk+ZOFK2vEsD67+dE0pE6M85IT2Z48RY
zJcpDY8z+UfLoyYvYKHeK6LPKU4br7Zhgy+JSzAbQcQEP6RL22wFoi0QppzbNArFy5o0HOFeHYXg
y8AVeNMHVHwVXOFZ4/9BB7fl/TS2MxUn3vfUyp6QguOalkoiRqgLeR2+lRbn5iWCJADaOfVwiciX
M/22XzK2BuoGdKDvyRUM1RGFBkVbkJfYPOlTLK7TDHXk9du3AryZp2wA+m7zSWip4SriLKwmz8DI
cyo61kPo+Tc0im9o0tfGn66jxxXFXPctMPx1YdQsoVv6hEPJkZxai0D7tvcAOdBX1m0RdltG1p4F
lv56bn0ln0crcoDxWYvvO8voAaMisQtbdglQ12zARGbf94OmkqZKTgKz5Tlgp99CUdMIJh3czl0G
xsnnVvdovoSGon7rjVKIPCTvXr/fzHCxTRx2HTDT+teAG6R8RkqNEuTxJkV9XrbLtEEm/TPWRyHp
FR8FdM8UudHc7Hqzbu3Q2C4mTIsYCzD3WFSZ7X4cweeUCh47f6R7duJKNtiUmg2xjthEOvr2Zsu0
SgljymcmlEwDJ8iYxtmyhxzPvxOHLYT9gMb2RMscASRTDMcb8MUAQT6KRBVMDdv+iC5g//qQJm58
e+ME3pD5A8bOAoj9keHq5YYd5X9mA98oYxbjs/4tW72BK5XiA8V9gwBL9noEkoYeU7pPZs5Q9cbO
HublTi7Eswin9JIc97o3hBnyUW1EnMx0RRoouEEwWCa9th4iM7aA+IomZ1lUM+peoFd8fNM7ScCy
JzcJxIlhb5C9wrp/UShvTmP8STu59vFENHdpy2qFfm/N2cisEVujo+BxGi8+eCbo3vprIHgK8992
0q9XyquK0RzyJ4/J4Z3fkv5lrdoc5hJAe2F6Rx4DeV4Cbjn+tpFEb/M9gCDGo9tl11wgIzGvbwwv
3UHpw0vdIiKSnV4xeXWQQAiqj/XSEAgnkxR5rbIGzzsqyGfgzvM8P0cSqqhx6mVoVyJ8ZjSuXrNt
AKPAXrdiuWtesh980tp73RxgculyVR6rG39ZSa9Hu/eyYHgVnPdC2ecqAXIxlLwGAGptVo+8KnFs
pq0HgwcAiqs3wC9B8ft3H+JO62xDmrteh6oIi7TD1Vm167WUvgYnoS4ronti/XD1YTworNY10xrR
d6Ek5l2AqbrQa2E91PiQGgoWpeiAE7rqrzeERrsxl7IA0KEz050+HsaLUQFb2t67E0Z6//kuScw8
U9BIs6ZIDgew5YD2YAqVzIsl7l4fDlt2rX96kYFQrdlQteLMikcUalvUfqgn6YwDCrq1M7bDDfwE
Uy8O/JdIFlQsIHNmlxCoWMMW2m0hHS1OThYS+ssu1U72gnAoU7i5w9GyBlIZ4M409XX9tQ6TXoS2
ZSDAceYDzVFlX+PwlEirL49DFXL3oydhCvFnDQoEAeW15dB0+944IWPE62XeE0GNlhLr3whe+DY4
0NQARXqLCEf94wF63IBJaV7Ez0LlWhEfgJsnfal4kGgGrEpjFNiXiXFFlQo5MX1avith3RwlfjCu
FxvD3vVI+5zYg2lFZDtmKh4Kwjspw6BMdeZefihD/p/2gtBJSUVGGx2lFRIxaR9ry1KUleF0ubv2
ROFyTqwv0kQ/anDIH18SN2FaVwQ7BiBoOC+hh7AzeRUAIe5Nr2mhEi0yw4CFdx5OAV3tIOJv+nXL
CpaJeFiAtlfWAUsOcNc6wuAe3ie/f3WG3TQHrSairGXSpF+q2J5xAFI4H+TYO6fxYKAV8fVMxDaz
7GD3BJX0UK03eSsVLAz/w29xF2i1yrQydzcPzY7hYb99Yu9FuZpHLMtVgD1lN7c7G8nsRiwa+o2O
30KH+51BZDp+vfFKLVBm3Hcg7xcpuEeBCOmeLcVqvKw4QqaZ9nHMey9m7lb0YoZfZbef+MJUoReQ
I8PzW+c+Qp8Ry83vJbB7JMHVHQyWEdLej31w4t3NS+++fYK8FRZ8IHEXghA7LGE0wGd7x8yBUVVL
ZQANTnANniao/oXgeMIJ2RZTSFTrOfzaBWEAFRQkl4C9QWyl8wJ7Bm0xhgGA1DNGqF9xvgIruJvM
xWnZvd0HbHNAfDmaa4JRUGaevvyGUZFoQQ0EiMNf9YaZR0f3uCAMXrxdCnxlx8Ef3USVS98odQWM
1DCVfknlzsB6vhaURF717YQzmZjlQzIdC26sz3M4BpcJCnXn9lbKeCWMs3rdAugYRJE65KgZevDr
BHxO3TT4QxN+Ngaf64aIO92O1N74Dk/jNxH7d2fpvwXrdGkTh9y7pyYdzunDQxAiENnhU0auZC/+
tgkdjzgGnP5FU5Lun3OnQq3CZRoXX2TJlzzQv02p18wvpdB31Mfv3WRl4cwIv/kVJ8mtbFxdQWc2
Fg8Oc1tzHb3ta4QY3ojf3GI5HytHcgFZxVhHat+63A2+mqSGUXYrC3aj+OATTDJa0e7LtknfAXOj
o7Wtl6TP7+IXTLSolEDn6eockovJwX4nWN9f3pwSY5Ww3Oz89OVAnmk17y36/ae2oAt7kMGTQrcO
9KimoImGULm6Wr915OjZapcOUJwPvhRoBxZsAW2CI8V49XuAun3m9U9BKEsFtA/PBdU88+iA26nf
CanGLx027EhJCd3Rnm7ezK4ddla7fk9bTrBUHdQgLLbyv8GDJb6kvLS8LESuKMM/280ubCfxFjxE
QYTGp5Sti7bXuWpsiGsqGkVSwY2NA4tUbuep3nRUGyQIgmiybX00E8Mnst4dhsT2dNc29pzzooPI
t3ytgyctKCYowo7RFBqvv2riFBq+LpjFAt8hTBdaOtmqeVHzwzcbMv/51c8VDHJUR+JCuweXseRY
cAS56UW/tXJsu21QdHDfCZNT3u2fz7pXNsR1+0G05wLDmCP8HHwtqx0v2iE/NCbZOuy1xNZLfntc
+ESeYR6OXYD8H8jqnKnzRNnyP/FVS2d/DpS6WRwOxtQx6HT79ai+NPAn8sJ1VfWAzHLsStJF3mBm
ETC/tPI4Vcb7WUKgOVsFv1UgIbLmriBgU8VafpjSZ6L37R0pkTwUHuwxYb6A9j8nsRP0fhqnMiZ7
7FnQtX/SpTF4zj0GJVdNVMDTFi2ho85ar5SrUufZAdHLcSICx0BfLTBE1WtTyaVO8AUcmg8zdJoU
aH7aT2QwLj01cDpfi9UtXM/u86meXOn3X0f5xh7Ec5yY+4twtWSMcKsUvQtZckcCQl18FCDeH6Ck
5WvFUTFHb0CydbdIQyd8ahKCiLgpzQ46J/4/uSNB1lSlU19LKZ7zow5OV7cEi/6Xdj9llMkchLbq
Q3CSzorcHsCNm7cAkvAKpEzFxYMKfGlyY8i0fve8ZAg2lTKHPYu3dmUcsupVMSMHqIwOEhGoIeHH
ndiXpubctClbYZJIZJBCZvyyIHY01umx9cxXSkFW93mdu7Ke6bGZ0lziAtAHasPj64KKUEEG2m7Z
IblZUjFj/Nxw/7hSTkuE5FV7vquqZZx9N8kASTuOF7H8CVLmyXHJFMk3deX3vSgNNSdGfKlKQcFv
4H4D+lY/pKUMSIG/bTTmoQkKKO6RnyGBLemZNRE20IgotvfhH43HVRulwjBonXZueCMdJncUVB/q
Kdps7Nd5lHXdK8MNlDKIPlQjJGw5MngbcMUmZOHrc8yGYZ+5tkwWZuaxQZRa47jcoMkpW3GxMcwz
OWe18sHdEa94wAeEH9/8UHp4NX92PKIO+3rzy2ivWBmyw86ZMcOBcUtuZA0b1QSDZXNv3rCGJ7XY
2fzd4uG9Ej0T6pLp4HdrI0vZcRfKW4+ZB8GWZgMv+EK+rVrK0rx+JUCXc+J/7fLqFmcGBBw3k7VI
vWIFI3XOZWgCGiOcKs/YDX1YwC9xwGaOE+50noGlrgd8o/MO6cjn/bCZiwSQJexuEM0vreV+h+dM
/mJ/W3DVQLgO65Ycb0jzFWc5dbJ9Q4uCDfSAH7NnLY2R3dXzDPn+B9n7nRhM3cjR+ScrK1wcB94I
syCbDgYUnwiBDcttZMlp+vH/aG1jl7i8PJKz0afIiZ4w9w709Z7qe7FYi+uAOea70RAVwtpJ/uKu
vRqFaJoNBt3cNLKDfpUzOeJ5CRdI3t89FUrOD+Kbjba+0iR+lMLP3u93kqLI8R6VptdL9G7erq29
e9QZeRXVSeCrxS4ivf8G57JWQECHus6Rn8fHnE+xs239Gse9yEaeKaGP/vDTAE+9bStGDVYR6T57
A6e19gLMGZXerJGMliWg1BYxqpIRwfzSrhUiKFVPPoSEf9PKKVMO513VCVcHT2I+DveCzlQYavlm
WKh797vzq2OM/nFDUq5ARMpeqv5o+d4Ej693Mc+Bp2hTCen7YhLLEE86dDm+wC17T1/Jv48HJn/n
MPLUi3fyx1kPP2rCDqGgIdVECl8cXaenHosouv5/adQDmvcYLVCHoKK7vz8ZYARxCNI6DX/25/ov
DMt41Dq6azPvTyuJVgFZFd2olNP33yzSdyvrZHeHuxDYpswZn7aS2QvcHmp0nkc8iDTzAwGqPcGy
m2KKiN6pOHpvC0PD6h1AcyRleRW9kVhEp05sdbPsJpJRp4EYPPAay79+mNID3genOWAdY7hao7gg
a3k4ujDlxVvKNTVqODVLMhsKrkDDomlKm5jLYNP23GNsHWFmOCPMkR6NFwDfhhA9zU7ybIaTHcwe
2vfAI1SWZpLFjyHIiKGjEF8w0Y4Uxc24e/Zrn/hLdmBYvWC+BSqJG9N4Y30sXz5BbG5mCK0Icki0
ZCPxwdoRK8NTigEk5fDwkL3nDv6R5oXNgcax9ceEBbmXd/7LAhq8z3FzTbubxXhaap76f18LgtOK
YhuImKym0yp4ib3E8CrhcIrefBMqWgdbv9lDtgd9Vrfj/IicOgwumnDFJAhDbl8ISNsaq23T5IM/
COPGjrx5qsoSWGdViaw7l9vu55exBmgyc8AtXhd8LTv5H34lGXbrum878rPM+w1izUtcJKdkM8H9
jaNYlJWOLCEZ2KcssXfFJpjJ1EiAeHpUhqoXx7B9+yKVZHrlLBjTmFPO6eCqZUtdmtQCLwHLyy9t
cG0IzAJoNt9+Ihc4nQQ7mZ9FJhzGu9bC8BQ41NbpyGWRXBF+zGIbA7bgKebJr6artQeMLeYDqDEZ
RQIf/6kqHj2lZpi7WqrDlGe2sGIxYqvQ0QlxzMxkpvT1i2dL5xZ4eRI7NENmlHtzNpN5QtzZfyKT
heohSEQooBZv1vyZOSmz/QHYEnfpMCfWXeVtkcekBHvfpMFDMf1wTC8TnPsl1wR7iCL5iWrHXd2Y
niDuYek9dINBmW7Fl6YCI2lAcHgA6hEh3ld6vmHiOGXFRD1MPfwZBn+iP4BtZhxMUb5oa4+/zuNi
joNV3CgUX+mskODUzBuDTMdCGLkNxlQCdUT3BnOMiF9RWMyf9UU9LenYQe6cRC2hn/1iyhaRpcKY
8dFlD/rIn4xR0vg9HwlZ97DTvOGpAYrE+U2zGtx1S3ttDQVi4lfMfjYmkhR1K456GvTo8HCuNMGk
nDVLqOVyCBihnJLhnWGM9Dbuc74UJtKfLBROZhCDIiURVIVZU4AsUlRc9anEEqhY+W2z7CnjsWIE
R5bW+sX8zEW2Jnjty+wAZwFatPQNcnRvkU3iaq9nGozsdSh/wn0uT38aIWtX4MdgLRoF68G9qytK
7DacFCQdZRUdWjy4MkYgpeHBD+xjWhEenZSMf+waAuxCI6sTvvL9ONnqtjIJDG4NnKbTcWWVcJ1s
62UjB2KbubIZmHBCf9s5Jkz6BhwyQKQU3rHxPeC9hLNeyP5LUZY8S9BCYVJ3J5R9L9/3M5SNSWQc
INrbG/JE2igX4Uo0h+N7kb8KaN2LXWBLVtATEbXgYG+x3Xe3gO9RLOT3nCP4A+S9FNgYElo00LeN
n+FRT3YD+vFEn9xbetkeebzHLkqwrVVPFgCmVLG7JOCSeD8YRr8K5ZBHXURuvJ2La+xbqL7nWtLL
eSqxxyaPj40VZAYterOF+UEJZ9ucXv5VPVc7+GbdgBxRwomx+ng5XHwMm99RAmur5FgffRgGHlPR
ybed+wU4brLE/h/1VFrUkoX/7Rg6VF174p5vlLLYuf/4xXUlIExjqeoEXt48z7qeIY8Zf1lIlCRi
uvcVRhEtqlLUzpHnihDgpycyl+IVJVh1UkRW2NKisBM0nJw0wufoYReN0TFRc9OEeeuTcNPR2tQV
N9gml3cykS19+tUZ6or563dANHb9h53hqhQpVMvItnORPoz5hqg6qjW2J7+Lz7mxOaMF1Tw87Lgz
J2uoKuUDSyzZ7Xdf7WjzN/ncIBxTE0sZtKjzpfleVjT8E8txwcPUsp/Aadr2tZ58w0sIW1t6XW1M
V20T3Wi9pESlRKyS2LRdTSdczJkIswTJkdq0XbXz8ysHKrGs+Laniq7/72ujwfD/evs6el8sbo09
MkpbpG0HU2FQ/NyUu64HD6k3k8T+uMgsCyu8B63uDIROyHKkG8NBpHesXY6loj2rynAmaFER/gJi
ZilBEU5FArbNWWV/Nul0g3LWXdfwsMe/q/Q0ZxvQ14ut9g3YIb3ZoE9tLTwL55Fjwsr0gMi3R2pG
EsGykukR83IjQZnFmEQJVIRaayoMRrwvnUp9++jJZcvciMYYGeqyxSmDbZ7xi3vuzLjMcPHlqJZK
z+938J5lsL5+t+9DuGz/r8ZmJQerTp6zkcpTAaclOZq2p+l461boT3xaBgmtpbTlb4DjpDiDMnAi
5qmW0IZ0Azl0xMWV6AfhVwHuCgcs9kAyddcSlZG4RzpcuTN7I5wFi09Yd2u6DNlABDAEYU0OnfMe
cqxNhaFH+QSrFC3UC/J+GpVFrtkWfdPzdFb0vpO+3+60jvNnDjS3YqdkmFbjAoJlT7paDRBoK4so
yTKwt9I8jOCwAemm91NWKoQnjCgriYpjKPgaaCfiQZSDHom8q/D7MTkEtasGfS0krhQn2rKUe6YV
BU4p3iEqtASLG9390bpQyWqRfAIBwQyj2Z2nXREjeEuckQ2ZbmVegFGy8rAx3kA3GV2ccDKOmncY
zuoh0d491sAb+5dY0wKUOEJWMDVitHYhI+l2taZ6N8uakuY+WXTgb1oSvb8MAo+zYXygH4RY2H+Z
TI+RgCvfufTSvR5bWiwheUL5XlX/6/89d3LUQlUwHYSlz50fIomTyntTlSSBtRwWSCmM2YacoEpb
Gpk1GfdnPNd9Y7j1X9gSyVozUoiC77Z4PgbGQuLetcbS/Zpin+gvKXu53C5kyy9Fc8CQhYvZD5Ef
6H/qeXh4pjGBorGI0ow/cXn2Dce2L6RtrBKNOjR5Xq9CsWXyZa1NpFw1ZDPpFf6ydUlv+enSZ/v7
Kz4vf5htgW5UqX0LGv4p+xpjD1TqoIgB+meyUy1dgexqUxwk2KuZWjodt/3fZ//ZMbDxBx9+IbWQ
B6jkEHKYXab3z5FiLSbU56cuFDt9oSOgw4qqxkthF/5oFOrariwbt+haDJG5wxtfk3gUHi/VALPR
hP00N7bBZjr+R6sgwxSprWvtgh1I12U9o+6YpAr2fBISR1NVtARqhb2O1sCoPQ1sY++bLPPYgP2x
s6PT1dRFs5HG20bo5B3YbUt2mswH8Sfhiq7vhXCzS+MhpASrGVtIWgmOYpzmQ47O67TjhgJNdre3
llc+5ALGDj2FtkPx3Vv4acY/biZi7WmQ9c0rFU91Gz9PCQNoZLTjy0GvMg5mdzkAx3d4hoxxbkJx
zzL0s/61mau1aJGWxN/NMsSzqGR84lpg4RkPm0JrthPVD6BG8TwG/XreOzJQQycAJFtknrahA8IE
0Vz/cVuxR8gbnIPFL6H5JlZHD+2Gi31I0f2uUdBpy5++XHLrfbT9DItT5YbtdguprefwodiJEHdO
j1PIRStaGCkgCz94YrDNO5PAsNHfGCOEq+i6lXOo+QA9J9euDswiLc6kIqDmapLy5DkdJMBjP7l7
POrpKTSU82ikmCX8tEEzN2eSxv0gP3YywsYBVx+KchhvGHVTnig2be865gH7bLuLVQRIj8E9AZ7o
RKIkRgp9F4RruoLQ2LsvM0/FN7SLwqM77V41lOox3dkAHTV7/z9/BPKp3ago6lSssneLXZyQeui8
h84VvkMtk0VGThAPmCp2s0x1mc0cUWwlM6hQ0hmgkiOvpVfBtUfU9PD1Tz1b0hevEHHTJ5eF+/T4
4ht4yPLxt85uEx3Sb8r2j/DtwcVJA/eU95+L6VfJHHhOH0/h/kkUNRpM48vu/bUsf3HBkHBr+MKr
eGUA160Z9vuOvLbjgq4d5Nwe+jdhJ1IO8CsMEq0ynqT5KvHIR7wGDJVU/PNyKbd6kB3am5GSpIHq
RQ8IacTlh1GdNl5FuvvUW1CDvVlHn8q8XRg1gMH1YsJTUaJwikfSn64bSk//npIcJLMWMNxHpCsK
P6+vxrV2Z4f2t2RbBw947Yi8mbjshDdO0VvAxtK2wQJtcy6X5NjOWp6pxNRkPAmD70fowz3/LJM8
ZQLBtttsi6+92ZdLXjbjfI499Y9W5DWXs479KUOWRqdh6U8G6dzk0F/WjeYQt6JTCfGM4enJKOWr
lQIDaVZCTTxfRYJyrT53Acrac0ULlr0when/OIn1t0aDqNSKeRxbpk5dP8YX62OIb/czuBCpsuUV
nZOygxCOyZju/rvj9+gwpeTMeUVAGukTp+ipBHnSEJslT/kQ97M5FS9/t3rtHIA/EUx3bwMl6sBM
Jn71Nc/g2xZITdzsuzN4feUdzFax4B+7i8vEHIisN/ZETQCg89GC0CLh+e1V9B+45HaRNnc02+eY
3BVEi8REk2wrR44ikegakeLDBoOGYt/z8QQD4GICSQFWZg8rp8b1IJpO2BV8ODOHQ54FvDuAx0Sm
/N4TvKMfxzpaqK7SZjfNetOsNz1jaxx4WSVokzLrGmyLXjdjTwTIHPVI785GyEq8F+Ou8VvXOaBn
tHSiKGIK9MsxjZpRqaHmV5ynDCr43u0cW79D1pXaZz17DK+osxFwz7Zty8FsPbkTjGhTuW6LzZod
0BIcvcUqwdU9b9+VmAEVLDTROCK21Xt7raNzqmbCfUfyjp/rc1p4s95J80/Bz103kqC1uglBK9WE
L6lrM+2iSHrPKJWoMmP9cT+7P7PoTvT6n0xAw5sLOpihSubg8FQBYJcnQVntS0L0sAweWQDMvoct
M7FRWJ2zmDpR2iHQZ0WixNlCVzoByBPw52vuJQvSPhfMgdEvdBeHLgkAsucYOjcT5PBc1RA2FCI2
rasD55m84LAtyRB1K5pcUWRoHDZYQ0Sf+5JoD6IzzzvX34wccJeYiiplvbA89hXQ1+UeELQ3phV+
PVinZirgEnnpO8qJDwQ0/bTi15wRSG4Hmft9NfcA2gmSodTNmmJ3+s7jVyABEMAuwmUxlwrDWiJh
V/nIverkWgi6OQT4FNg01i8E8Vaqx0bdPC9VJpa20mTQSdeOUc0SDq2/D48h97ziteN/8nHyVbGB
HVbJeBwsXqKuOvqba5PVB0nvh++EN9dWBeg5HHcD6fGhbXB/QgRhRgRGROBZ/WFRW2G9IRV/zf5y
HN0uQQhqkqCCyJbxsBEApf5UTe83ILzFIcZMqr83nuDdYOFndBWShm+UVqp+DOG0x6mvZgOi9goS
xT2DO/NkpvlrpsQzFneQzr0QbficLdQpIAz7W7XJT9B1TCdPbQNECL4uRQhyVscz1TY+gsfkwirZ
cQBXoIT97ZFPe4mMqRp/Gjn0BPgDv/zEguFW89NV9BlGZdONJPKFY/WLnUbzGDESDTnNa99ovd7C
mhLYg612BuB8i3ctEqHxM5203nzT9g0uFzFjR/MIz0UabjqomJRGm9swCplON6eRcDGYse1GTOeN
Zb4n6gehMOce8nIj1iVktPAmTOtC2H2P66JeUV+Hp/xpzLU/jwZXGft9tFu06XnURtAxPeW9zOeF
RpWkckUAKgSs6/y4aFTLwZHaodjFHuYt9aMcQR4VC58s1F9lirf7QHLvzao9qPSNNJTc6RpsXLHx
g3O6J1bi8qL8ZaHTVcZHB5kbLUUwHNn7aEJHe0MNFfaNqCaOEHzeCHRROZyl7zKGI+dX0ZgxoXuZ
TITfl57b81Mw/uYxzx7YySTLMg7+nzTCzkVRqh9E+hAwTY7Z9QOM3+v56BdYN2WIQslz/YMNtvjx
gK/se1zjngiN41IswryEITJDs3h0dbF+7zl3fwCleCHJbBfsygTnRfinE9zz+4wQ5XohlGkw3F9g
bvOOsuZddZoWtypjx1EM9j4nV1I5dqHyafQCmQ7k83CSlJxgijVImvRRE1VDdfAlSOlXnjQwN4Wy
2UBQ4sZNfOYB9nIl4XITvU3FHcRDoSpI2xt1j0l48DDI3C/COVhorVn7okUNBKflYQjbwYEHpvcP
560ckxwr4LlDVUWfKqh+AOk8ZlBKGidXqlOEmWUCMgG2vt6O4QDkaVfbWCxBm+YTQbje2p8Xu9KF
ptQ6p5ajM/WdOW7gwermETNM50F3d36U4RnxgdTj4IKUYAm3aGFiXqf0Rr7d8iJONwhTqKif0su0
K3u6RmciVOkyL65CQDFD41lUcqv/rdDJP104DUliofidCRNd2cfwTY3T1u2mC+g4mR3dIbii0k6O
ptGqEGDnNm3mO7vWkGZg/rWZKdXjYf9VOqLx8GMc4GnDF5P1xZ9WmeUp5vzBMAPD5e36iIeZCBcG
/0i0UO03MUxenCfBWbGwUAzEKxYaAmTnGgakAHaIApierfDnA5Ts29P++xLcm8QBzQIkjUPKqDMB
Aqnk9dkWp0hUneqBjqBIt5wIDwmJV9fnIH8z6dP5EYdhWFH9KG4zddnGFAc7ST3Y+/un8o9biuvk
/Tg9gt6Y24qs0WCM01ETdrBaCH0JEq/PJgnTtobK38O5wYl0xhWAlFRvpKJR0+h5f4w5TVmj81WQ
+p5bUnf7UU/r23atz+eGXigVNW8DMJeX0SOqSjtWeWbF/fzpKP35sw5e/xIzaAPI5qr6h9v/iSoV
pahQwa2OEUkTJfI3NoSkJoCia9/7TWCHBlR9cYoPVDHP76EBt0RWzLu6u7859MfQxwwbwAOTOe2L
kZ6OSjpMx+bknimOZhCy/2nEzqKZoOe2MyNPdT+Q5CmH4UcfXwxk9yvyYBJ3IeQ3GJaqCvj4gulm
wodSl0WixjCeOwqyRYvOMoHPTmCX4zynZfZGkVE1X8clOUvltpSaoWsDXIzzSwGom5UdsOiseuZI
dK0vphG/QglxfRRrf2J8UCjbl5cg9nfR2kY4CAAagw1ZyMCLPXMywOD8ynOtmBaKpvcDZIRphDX8
AZgACHTUGrrC14GtJho5xvwW4dk+AMBxJgUAS1uENUc23EZnb3ta4lc14tz586YMyyuwveEJDIBI
lm6MqBfz2ki9IhCwyVhlgsa/r4WcsVDGSsvZyhejJCSWWE8UoID2FSJJp94u3LxM4vjZxD8pWMCc
OwOrdvjEDGtDnG6ziWG+LluqXkJ9Jry/qm4YyR+a8UkTbPZRhIg8pjkyZ06EVxSVPUPKZgDOiFRT
gCZ4VlcEZQkx8L1iv2ayghXjYQUY44OsD9fbGSMUlcuHpvgucqhEjYMUdAHL1Ypwm2eCgdEgMTyO
XFhbn/Df1WWLhOZT+NUF133TmhT9V48NyGsibOtFIeSF15XgYpqECuENpaFQb1e6xZf7iL8R+J1a
T9I3cF56mKylk3OU3OmP3+w3yFlQgP4kORsoc/lFDs9MxbOUBR86hsBuKCGhhrTy42Qp4y5k9h62
WfBbL1yDoblMH/8PX8S8GPtzFrnu6iMT9McFqjxITQdECc56DjOLX1HYK6YX+jOhOHPliz1PYoCX
4CUjMr7pKTPdj1g+QOMy9vYRb8HW0Nhzzvrn1FjtCvV8lIjQGlm7MjooDNftyFeEOQWVqaMJEksJ
OoGrpfX4YnjZIRPzUpjVuuNKm892a60G6vDdnLKkE/M/k7O4FVxDIpuieGXKnvWFVEBk13eE3VNI
nzZVdaKD8GjwNXUfQ/jh3PaKOWPtw0MJ3JcApKA1DYFWEa7THOgNO67zxIxjGOzyLyRapRSEh/V7
m4vR1DLNPeMAl6JMecn5tEAMvnalHFks+dlssvo+za9YsmUXQBc8Ib6V5UxnRZ12sJ05PLvHDYZK
P0T7pw/vTZs5gIBggjCIwPocuvv8DyeedFvLTUQ4Fon2riAxHPsncLlT1FwJdZ1HyiwQhSJ0YBEg
sFkajk+rf6ZZ40Ie6ej00dkFv615wh5uBqQwcF1Dhv2huuG55LNAYuH01EAECcdOj+tP3er22EV+
eaBetXglQNm1ud8JXYl9ecTmHYLuwAqsklM1YCuTyEqZx3zvDqB+/5A/YAoPwxdFbUaTLzJTANQU
8nlGcJvY7JHD+SScKWUUozecraVxF1QU7e0kbgNuzCviUXlv6LLwYUNPOrlTw547iyzFklYbUwZ3
nxF1oQJeMjES/lhWAqBdhheTMl3YWdsWLH5060zpMhpkIHMZoN+EFDBDovIx58jzsj+Zsajk7rzU
pusEafSO21W+i/M9VXJj1Favro25gFs6BwDY2zFLmAt5hpaJsnEnvOTSB5xJC1UjfTkmIqHokn1j
a3XKF09ujalOB9YaTBJEKmeGw/CU7KZzDY7UTVRbm88WKK6LmJ7xjJMt+CgBDwaDmah6hE4fHyJZ
un02u97IWaCt2pHwG6Ls0uZyMeX1RSmHR7TPA690a0fK/mc6oAEb8x2szn6PjQBW9WiC1vaSS55l
BSUaWzZC0fuR2Ih+ArQ90erJrRXFiHB7ePhW1JbYa5QgyT6gdSlEarqo1EuASO4MAY8opIilXWk7
pV6cGDuw1mndZSXQIPblws+Wh6bba3GCu+L8cyNwISoguz3LAdX9AKS8vEh1DhkwgS0JR8DEfsAh
X3IQqnxZpjK3pqE7EM7L7i5LXWwtk3Kyynk/BJuDwpCk+a7O0L1JAEqyHzXONj8/+RlnUzQJgLDv
k6VRTueVM2RlXE/bv5QBxXHN9eAnnVtlwWQ9OBO2aNsU0tpEVmb4muO4REX019qx42+RAVURF2pA
6UBFxVfMpGYENdy1Wiqy6p97vGkWYSmMDbO8TH8Bnvkc7km87B0fJypstqYkEQmDjpNYHOvj8hWP
9dtbL5qO4MJdMmuFp/FJr915TWaqL4scfPYjL4bpbIxB5X+lJrVFL2/hjqhAXe2bEUxN7QDtw4bW
2ncfk/nwwTKSQltKm+wgYL4xQBNO+YMAplhNSa9PuNrXcraHS4J7H0z+v2APJqTbxnodWsAN9l/T
3n6w3oMX9wMp49I4Ff6G1wo47kFuB13eHr4/NElWst1rfwGg/AfnUyHrBw+myFoO+cogyo8cHkGV
Q7ZUaoYR8pEkIow1ejLBQ6maiJVvMw2PHvypHcGhzqsO/wUHx3DFos6cIIA4i9Wm9xBxgpGkKFSw
XpSNwMcP/taTttmtf17i55DlYdPnryZmQJMJktdje6UfK1anyNnKxvqjB9L6hFHeLdIUQHOlT1xD
3AZe0h+Mdr27cClzL23cZsRu/vn3FNpES15XNKlCRiBVe1qcRLPjQqk2NZU9l2y/HZQ1YOgu573m
kF3UonowGNBkAzI2XcttVCJlpEcY+MemieJOqrT1RsQaTffvKEhJdY+4J+6sjzXe33Hva4RsfU3W
oxI45ktpkoLsux9TeXsGv/naT7pq7qFaH1Q6Fto+fQBYQg7/QslPsqtbYpzqDchWbbfN8kZHac/y
61NEsuaQPEpG5oFdEzfdveNfLCJLDCkRii9H0KLKvbe6u9mQuQEofJMkkfu0Uonm5aaazDhZyE5F
YYWirKSx7uDwQqeeiWVZwIaSSEYDt7n6V1j0x8BitNIAebkrRaW9ArXJZ9UG7e8ZCKGlxFk4YXcW
/S3UFZQ8vc8Zuedgp/FRW22wEE2bJzCdPATZuhZ5Yptp0MgtxYCs1yZf7hUmx7j0Ict2ZyGeC7Qv
U9SFyN703zNM3bdagO3oc9YiDd45IOizbY5V+HRYvVLgoN/Ae6g36S5mrHX75RC31iItHSYmmQwi
B0COXuE/wxE8GZI2jvH9NPc+KtNcrixJeKPctxcbcbusr0IACk9qKMhV0MiMfO2OHDeBS+MZVmso
WakArth0k6mZNhOsuGvApHen8c7/yk9eAAHTgUdsgb0qQ3JH/x50O9Ubp/MBnmelcT+iLcNKJZek
7HmYmYUO+9wWCmsi6ouX51iqmw3Wi6fywPhXqSvQcPUrkRJIcvFtGWUmNgIBgXLuJSmf3sPDsWxv
oUvjhlDFsM1+hYSf56gW4ps9L9hvTCRfUlr/vwwPH9rrmv5Hr+P0cI5k11K6tqY8BrIM9zcR45bM
rrlZ9jMvm7Th0SEMpWFVc5PkTJR1cgnDW8nR3s4rd1OV0V0SrNFreS15zGxnDxMFhMDFZ6FsLn4J
GehfCpDjXAMKdVqmGmI9llwR6WvK5AKVB0o/wmDhvqZaxmqMRDgKYgcv0Q4McHammCgF5QyLBqKr
ADqN44qg6AenLRWvlcvzyBwJcvTFZYsij4dg1ZWA+HfzR9e6k/kzJRg7OMNrG3reYmo+au/aXapl
W9BNvvLWu7dZEsOQtU0pcgeiRf++a1qRJ7CDbipVEAoEziEBWoSIKBQvYD1WUdBe7K6RUmtYtvaC
UnsvK4KvGmZI50Aho7Dnw0m0oNKjWgWu/6azTlKJ1TUlIXm85sLljqZ/izAC89ih/DnsGyp/P0P5
5YZOB6tE+55HOTeKemQfZZ08ErA1fFWuHGEZOStS3lDtxOfhiimn5tUSA8pQAqEvoItRY+zdslMA
H8u4F+2Yl3A3DeiWwYvmwP2v1bBojkwht3hfzYuRDosDjQ38q3F6sVTOCX3cZuLot/nJfIMxEzQw
jETsvXqAmPoBWEZexH2yoeSK7PV9lfLE3KW/PpJk+ja9z1ATv6SCWtZupT/QcZILc9ai+dPDWo8Y
xYHZwmyqtXFqElqKtyOu7XULmOMT0xvTAWqmmdOoMND3sXtoyXZuXJubEc+4GSC0euSi0EBGj75l
NvrY0kzFvmBL5jaHyjvWz8lMjbkajP5FubpsHuzpeQ/9s5IVKRZbPBMSkerTmcVIrX/RtD1mn1st
rhR6VH6MpK0X9u/B6O975wc88K3tZKl9Q8xm18VL1mo+5zhDj3Kzo35jaJwqufmAnjH45rHPIoS4
YQ42RDXiXgziqh00E2OBjIlv8BPok6ZD7mcC4PiLVEux3uHywzNM3/6XsO2pr/rdBWiC+crjPw3D
nDpSgUXf/dZUvaBO6A5Va5fKZGJbwXxHuZGaX0KpOm2yNGwMz/Ad8CodzNWxY4SSGYnCRwKcg1AM
lw+4srg9pdCY80iXrR8TOsGKupYDYSX6pCnFTT0YjbjByBQ1bYeHwdPdePlVoDbGvkJVeq/o3J5F
0bRFFWEY9C0eQ9Iq79iQrFGOciXUkUPcC0kUUrnejeuM5zybKHILUCToAnd9baeCzFaGvN1b0zdC
taGME8A6dyAnv+5RU/Jh3fKBUc9+MO13k8qnuhHQuY+5gdHxkAV7Ll89SwM8RC7NWbzKcRrfLn3g
RDsD7IMEEBFd3WwIMPX2MRTZMWm365T2jLpUiAS4/Xqy94WpIvdUjpfB6LgvIhIEmGh5pLF3CENZ
pB1b2M8hEQC2vR2kb0luL4V4xYGsYWkepCxGmDeSHHHNPZpGl/di4YwLvAlsbRiC6BdemR0v+Sbb
LCDE0La4p19YCUqG937g/2a8CgBaVVAljfkXTogh1ruEQ/JnNCxAMkAfRU3qkugS+uUitbiBYuqe
7lhovNQVGTyLvcTsO/X8XGRjp/szKgsIV2yEKt5t8mJKRQfg9ACRIjjjvcl6D3XKHQd11LcF1QsE
GqbaChWjKx666z2pAJL6++nPvXQeFkzCFbnTDs+2xf7IfrnV7whJTkL416hcIZjtiDtwc9Q0Pq1x
zjr0PMBBTfsmPZud+xn58hgl+9uH02YSMMQu2YRZ3GFS02/mfOu6QvKH2vPZ46Bn1m5IB6G2yoaK
WGYa40xVo/MYBNvW0Krlg52O5ZTIhypfpbGgBZf8uXbvDYLPWq/iH8aV8sAe+8EyY/thprb1BzEt
DJljx/G5f9GJ3cWcsXq3QC6JmeEtk+yhR1XcWCtg8K8LZCduAJ6DA5DdcrRQLqm2ZYvIbzktQdob
F7Qo3lROMFQP9hAkc2dbPbB9JbBJ4wgHNxV2vF3ObOiyOg/OJRc1e6WG9Wb7V4B1A5gS4gYgAN3E
86wXfXq6YTUHBgFBnsmtGDsF8QeHTlBRvqoIsucdhDwX/xOTklZgQhdEjdk+PNOPP49q4Ivrnk/G
cx1kGrFqIS96s/7b4mh/GA6toVf5NFDmBeBbaotXkXHcDAtPhVmTXLDx6z7GR9tvFnMZZm7+NaXg
6dAuwRZZd0H1o9UA2h+neVO1QHHfvAFR//gYXE/tYkcbkvuDSLgXVxbC+s9F0x4XUNYTSL3IkYXI
tgr8HQR8ClYLeyK0xuhFusS0JxyircE2U/yeUbLQNAH4DVIBOTrJ/+4QrbqkAbkF7C5ryJjX3jHO
yduve5kWp/YeMYyLk2aepi3wi+WIlM8roluM3XpHzAlOp7gqYZhhrSEa4fd9ijX/is5oj0TDx+C6
o+zkuxZHXBm6gG3AbEJjir/Vh01ZAETpbKIftMZFT3GaVdu1+BmRpDkaWLPHiBnIvvklDwjRyJyJ
1Suotr9TjHSxgKoAy3Yc3Tt2qUCoQ7IErmlyRlLqQ0E7QCojJ6a3db028xSzPvIIeuMOMBTGcLp1
JrAZiZgihzlkFI8MA0KbaC+UtVrQNKIaXuGqfOlR5JIhTrvRVTx3iCggSVt6Xomw3UUrs4Y1h2KV
ZDLN6Ai7XetiIlNdaigNkp4UGfi15uXiAqhC4vG4XXAJSb6RTvHWMDbiLKiTN3PjpJPF9x8hq89y
87cShojN8QXMDB+oNHYDEi0hJSJdMlKrS+i04hLicRjF/uTYgfLVvQysd94gv2qCTZ2luusN8nSe
xt6z2llg2BOHJ8tp1zuWD4MJPx10aQ/GoBqU6KUUK/HhFBaPoFG1rxzvzwHRX/qyvQ6Y90Pi/z2z
kchLc/xChkKTh1pFrJKU7MlOxWXZ7x3EAHQJyaxqQAOpzMrmnBVkH/syYdMnqeV3ae+lU5ypkua7
5EZkNfpDvdwKJ9dwGHS0T12EPciQIGcLlDzTXtupvXvDRzvCejQL40FEYYpyqLfZoDYawjwfxzdQ
oghOnY40r+C+vtxnzJsYMQvoLY1N2mTU0HeGDpOpNQ2HEMAlVu0EmhzfExNeu3Om6+Fc+Xy/a+Oi
0OmtiYJ8qILV8YvQ650cGS60nXZu2bGtTYkHP1ywPvATsK7LV3Nx4zChi+lL+d/cLUPXot3wuuQN
fCR9g9HYogbpqngEV9BAZfljzYxGSC+poXN7OJLjBjJ8cukJatr5720wMFXbgK2Kas4BvVrngeHh
1lcp145LVSrzlBSe+P4xuiyabyJZsXq1PxQUIAadWd9PvkaKnNSNQd1SzhY9NnVJofu5kT0XQODB
zMK5jRLZsaAtKIVbLobb/755Kt6Z8C2TV/FqO4t+TBBOcFXpJ83VTT6nZ0ULU8O9wAAnYaKAWrV3
6JSk3ceZ6VCiLQatJpJXKE84+lFNp2hFQn6KrMYVpG/u818t3W0JrwOL93OATaOprqd0DLncb9be
Wi8ne5y3DmGM94cXBc5zU4PYeXJEU3J4rAEoPuzvT4Nb+PSBQBnP+4CpzJtUtpn68Vpc9kxwRGbg
pZ6QRs88cbf32ufk20p9DoPI/mONZtHypLtWxoqvZrNWML4aFd6OrFBePJwYhkECslchRhtUSxcu
gix3mIFGtrAGEjSNLHVSbdiLubYqy3D9qh4XMRVNwiqUnk6OlBah9bbaEPe4b0DDrcKSTK+zlw3u
ujQfWUMxYAXs5W7B5aBwLxEMZgz5kx+N1CwlrQkZRfU3kyQg1P5d7/kjeu8FKw64AM67KoAXvLrD
kne5KtnarVxtU3f1EA4V6eeEtiSpFJpPC2iUCE92K1yjD0ciIOEd0/2g5S3O1EN19bNnQ/cHtzNa
EvbYkEeirO1kU/Z+RrnsPIEdMiCEbhCxSAcdQSuWX+DKmYEVZWcOh/xmkDKBQCCIGEI4JGRQ4PlR
HWcIH0JxJpr5DfP+hjU+5oXo7mVZzN0c/O7cad/40i/4gLSnSNf2sKJVpISg+q+Im7ezkmgucBW3
Ow5y8a9i+Ef7qI1FCmeXgGygXj0GiocoFkBQ0FaX7YcXS6ZT7yq1Cez79cmnE2pFciqtbC9ubhIV
cvc/Th8v+r/fhJRszwAz46CVCH00gMLSDGix7gQSLm12/ifvqa29voxKXnkB9M5e1YrYtOn+u/eW
hQk318wvekZUBqLfmIEyhsK98YyF6jL4SDScrShrXO5Pc7lxQ/uU77mdPvmsm7ckfD1HpwevDqG9
WCSxkMIZl7NUeiSh/5rFgs4QvHUNdFnvwUFSjURR1oTsbvArtynThp/9TCfG8/D5p4wp+tRoZgxC
JtfGHTc390SAlYID0Tkyxd3BRwH0qBce7iUGkwW990VHgOLPCgZsGdlE63DN16onzmZGZf1PBP8v
VcdJfuC3m6yhwO0afQaID38I4/U+qlBTMtGNPR9oeB2xgYY9rNQHdqevvkcLeCeOK37kS5m3hvpV
YHFRNZKqFal9tDoOSSMFx7OuzLWs+lzhMH/Hb6z39ye/UXjnhoD3fVauPCsgyM5GddR4hxbc3IAy
+V0BFYQsSsg2YZQV/v1MEoS0oHbP3oWI7HwZsc1IYRIpCot0q5AkMI9rvWaFptDdUYEm3HFYgr63
drK88s4w3lioJpAlIbVSw4lkMjta7H+vQYf91j6hSA5DLLivk9XtvN4veUCVyKMArGp6pVSbuPap
vnbF0aZd1+O3QMYwXNgWZdTFBOieVvP35Up/C0TDNxl7TQIqQ0+xNo50RRkyrjkLZL8iij9J/IzS
O37mlwAd7BA13tzo/l6Knb6aW/rDB+nfQMgJx7XaTsidjQYfz78yATWJHJzTn83A9KJe7KtARPeL
fFmVZrwVy+mg6GdJS5J7oKeYGcWU2W0og4xbz0hUG7I/Nq7l2h/RtU1+gkchehPwAD8xLhgT2LnR
z+Q7WhLnQgxtZIsCxKlilVyXO8Rrya6zkt828AIFl1fGXRbpcHMjT0KGbYFBZneq3aBZRFfhP6D7
PJfFy7jIDHDuVxvfMJfpPqtuf/buSKrLW/JvlPpKecU4vlOajmGDD1vdczCNpq4LRMGBp+RW/Att
9fvMNxpi5MIs/K1pSoFhpgueutSGS9pznuZEt1SrUv+1XrrstVLzwdZZM1b8r+Nl5eSAcMSG7hCl
W7Fvq2muhawrOdF+ACcvHwmDqFLVp2HjyNfL2E9mNeBH8+FzUfNq5BixkyJgmkXvVaGYjY3y8Lq1
a/1IQYzdCFAR7ZzN+xb+VZ1WpoQ9LsyVP0CpLO7P88bg/uYtnUOr1JzaYOuGKIjUXHQ3cBVSwgYx
WuVngPbOXpQ0KPL88ZVz0oaFORE5NmiANWqhfvSaG3rGq4ej1hEyn+UgQzvHzFEIRyiwaxCOR5j2
xpJHcgoWW8WSu1Zvop1sTRmh6bOeEy3f0TBzKClMuNwV77Xx74uHC2Y6lWGNDsbIRjnwUWDVQKhx
efA6SDyTpBbgVuCjBMkR3YHQ69hvQjeZ1UkImyA5F3DEicAOCbkuOw0Dq6ZcxMvNiV0w77nzy3T0
pC0MMz6j/fv5hut8Cjz5LZJPVTnTMr19Ea2ot+hELXmP9nXX1IS9KSwaB9dQ2iAuhEVoprOwupVL
cCRDDSgFzrtvfzZbPLhIyh6JY6ddIROldCrE8WX/dpkmQfq44XXqcCVKMvku8Bfa2Zw8tYdw7Q0F
3+R/p5q4GIpKN8UFR+GGWWgCyupj0DhUHtlyg7v+X61OOX6fcB6+lFE/328phY4MzZX/9zfl9KgD
RmSalVvPizfElYmgRMyvo9wxwb9g4DPHIuvny0QQLKwW9ZCurG6bwz65jkZQdGkfI/F08hmg+2EM
dr/siVJaWP0VUkocnNpN7whafXkI5IXmFzp1BZ2FD9i3K0Vjo6Q/OXX7D5VjHZ4XZa6HWqgJFQ9e
ewQ7uvRAoC66e6TuVB7dwR35lpzMf1nn19TTKJ6kMs+VBG2JZ3ZWvujT9iaokAEW2z0RkIgJYNlR
jpaOZzPurZXVeU3R7XwIxIqwH9II7ng1RLp3nnrWbgCSgj3FFpaw7rBGNNNWxLWrDd3lNemcdZv5
aQz98G5kHnJR/3mW1LAaDZJPQNEBYkW0Rd4p7zviiPQlBjHWgFSnz9ih7tcq7YH8NHFNamaCJfhu
BythBAG4Vgo53kM0SmZZmT4BQsNpMim/wvEM1b+O1yyQlEEMPGjbR2WdO/cSd3YddqPn30l//ceL
DO36PfqZ0AZsdH37m7gGWVBzKKx2wh/xeipCA+/H/1d7bPjfinPFzr/ijQVndaRSe3iLww86mfCw
6rhLd3PA+bSqFMM6EFhiLYYVQTDA2WN5ZvpU3AhSp1zrBYiYqxW7UTwPrpY7xOhIAoPZk6W7hZkc
RKJ6hGGcaXDDMPE608ossc2DP33qB3lQNHJ7vVOL2XoK9SpZdABmY6DN4p2RhPscQiC2JXb4hSv+
488b98MMV4DTzCxxVr+Pym5I16E6OgNkDDrNAWEJieCpuWd44pUE6c7b7ViwmKQhSL/g6rDRCNb2
KXKiggWoAZYsTEYOM5k2/woKpghhrPf0+rdtGqhVcJ9G0dr8cWWMqnEcuYpAWnBo5vvm3mUr0K9t
SNHleEyeHcZKxrsPYwKwiS4azooTu7R8NCagOk4sBgNUyRGsrcdjkLAA9o496di6QFezOb7Iwb3l
mJiEvILZM2MvOO1rDxqZFqQZm7XXxxHzb/LSlaUWHzMSCfmkWGkWinXh6GbpjN3rNU1ES0uvbiKE
q7LoEFeEjBXd3bpoIYDGfB7C0ZyU9rH2xurXIQoTr8XeWIgyONyXWzHlb+Wq8JUUk3ukW5zjFRLp
t2x7T9hYS20Q03FtreQ2Q+/emCmD9srtLLOhrXIDDCyeppmAI2gwO+2DDkISkHd7xJWFbohqEjl0
Lp39zHNocCNteqYCeJnFfouNpvf8OY1dCTp0Qpjv5aVh2ntWE3KSCuAc5CwDj2PL4/UDYuEIcW8i
WNAcLcLLrTjb9YhY5B5XxgO2fT/Sthpq2zdILwwZ/Wtenft4NLNuGxR+TsuliVenZjuF+vtALiJE
0ur6sIZLD7Ofke5gROWBB7aOH+WCnecexLHeQ0wXbV+m5fxA2q8J5nU0lUSQIkuRnM6waEPlmY8m
8YNmuRheXnvbilEgzZ7mrONH7pRVQWZZLhmSxWrovxk8y6LFYKMCbsbMw4m+sCBO8oNz5LrcODG2
pJa+kudcCRa9jt1DR6iL2x8fVO7+yQpdAfDvovcDQGGvo7esYc1nAujbqzTyshYIjRs5M1vunQwb
gXm2lqj4l5Gqh4pQ2SSiuqus9HAey4A5+90J+LbGv8Cpxv6jB2Bo3CYp2C4pvXlh3hQr7QwA3xsQ
TWal3TnIe9wqDvq1d3NelMSqKhFQhozM/Rzgn88e+Q2uRxP0Q6rAHRwtfMn3ryMDjebG6YCq0Zpw
4M7o/HcodI60v0nCjhyUwbsw/50tpOFOQ1LFxnObMYqfg+cS9KHo7CXG3FtKD7k79G9Cnt9czPc5
8bP+UzUZLiXw+xUiBzPcxrSe3EFfB9sAymufJTmCIzQBGEFsvK6u/Vy9SOFLxRSJ+KOZuXCK+PpA
8mKPZUq7vYexIfPKtTxgS4PrgcEZXaaBtW4+GNzz3IAlILJZvhnRDbIu3UAuP/9GoNfbk7PpM/ni
Y72BEgzs6PgJ2gS7Evr6b3sov573OICsLDnXIFVYmGKHnLWpJ3oafRhbN+0JF8RsXEqhWsBAZXvF
sqiftjbtFDOoQS55qphMQ5G5WNYjVc/CU6RWmSrvAx3ikZVTOHpBhBHq5K06Qr57KMEU1ww796h9
awvQyZ0zb8QewNnensZ7nfJuAXLpEuUKqH19svvq/TRyIOH6ann0tf2RvTVq/zEYqKjlOeRvD/ST
ql3p3QvLNpV++WYMSo/X//vyzX5kchFQ72g3soiUyX4PYPHUGzKGcvaLxvsBgxFzCkUbfUDnDFBb
2WK9jPz5Oaud3N9xucbvfsNnQHUudEmWNkfG7SsLlFHdfhaDfZ0/PQaliXVitdyosTVBqkg2dkgR
Rl1O31+N9g7Kk6mcyo1m59BL5yucx2vS/ahsnWVEcq/fjey7XkgCWjl+LhSj+cD0fwXUNu+dXfph
51YzlT/+FRurwiTEVi5Zu4o57B558qipxLHQwpzj1ON0etz5cEi5gvFAeqMNU8JUblmfemTZKg1a
PFvXztI/X9GrSa7M0aufhgpykjLsHqeyELN8wzuoEtU5yk5b6a6k7Q88WoHYYgLEm/3OasWrAgoa
kXugR8J2zS5sBWQ4VFAPDWe99g0jSDyQJrM+UImIoAKSJS0sCm6BWDh8nbUH1pvhC4dpAGEPrYtI
H18a4IumPrMncuaLsih3uW5xrmf5hEbXU6defth0t8GGA3iei1mXJbUeeUzlTZoG61SCgyhMbzTk
uyTtbTiELKUSJEicVRQIMRKE3EFiuGcwENYWFPXJ4RYVU8wC3Vl9zXtbfXORdy//p9gH+A1A2wXH
4v7CJv3r85vQGQLfB4ZhOlGrMMxdtHF5+VIZAMUfkRM+z61Dgeaiz/iXwEkF7XiC4jQxSpaB3pEZ
YAccoa3ifMcnbnQum11JusEOXeQrVP1MViyB8p4C7SiHWDTSeixaueFlwv3R4V1t++ugztjlsD1t
eWLorR2lGD0sSuF4Oy4OIAHE9zVLTCGcvrnRmUmmAlZkpOlikF/zML7u/yfsmlSNte1pS3OgqPmE
zj0GPUzxsQ/HmkqeT0rVLCUzGNBOCru7vW1lfN67wxvkj1Vp5m53DjqE+j/zkhfMwYm/+xMlId5f
ENTkMs8k+yNMuRnQFr+xdnRtJAo8tPnOCqBszCBSUJHx9QLt2HcasMekMJIynJswvnBlMpAQvJQL
z5d3AlXLPV/w+3sPBEOaJoaFXBDUrrSMr6kwmoWLYt3xAClANHlepABja2i/SfxRbBMsArRtfCLF
OSVX7n9wyYYb1cQ9QBLQMOLeQv455QFklCAXViRZHIAkuy9ffaKwR2VyHS1oreSEc029rlyCKwJA
bnxi6YUxKMfjAnJklB81qezo9ENpu9/tj+IguKo38OnHoGFEykRuh0ZPm2Qn+E/jgFTYtOinCvF0
wlF3LkuK+mL4EggR8OoYDTamf+q7W0nH0QJUE22creemt7lftSPyPEsubFPAUuS9CJ+hI/2TDS6M
WSf9VX4aSyoHXxmPq5RPZUaL50go2hFNEEQYZ0JzqgHhoc0qwOaOv/ObRED1JFcb2x0C+qU/lvnv
FZugWZFtc0n5MMVubJuWNEaPdFoYcVBrQhUCcM6lFIz1vedo0BhaPkB3tbJ91WDcWGMJY0H4iF2J
qMTweuWMSvyyo6zHacUuPtn0vnH7d16mZvEOhYYMNsijn5GbZXNAAUz9pNMkWKe6e4i17C2Z+eac
QT2rhPi+wrltgHU5pvHTaAOgl8JgoHymMSnt+0HGLQyHPw0vvClcRZ1eW1YtvUnUB71bjR852OMo
HZzWriDjk11hRWPoihOlxfwfd327wocC3vGzfSrTc9sE51W1mbf14WL54Wr1KhyBW2L1NAYXvghI
zRNwpb6riIMJBSDdA1hX6/nF6xuhcOXeG/OFJgoxlrOZzdrK3uw8CcUQqs5gWxTdGuZ5UYpCX8G7
CDAWI/ydpHvWMV6fBk7xHNs1vmYZkCT29eyLANTVjNQCOheCV1QOwIfICbkViBRK9ux0DLee2txz
Gr93/46tgVR6bqL0A+6s39TCWsBuXTtJ0bqPFulvNEZ2o4FUkEiNWD2X0JXgQ8zbpfOPEcT3S4h5
yX7/hc0iB5mH0lD6gQ8TddHGNnp8OeCJ2nMVJU7Xn3vv0ai83yUIm5Qz7f/p8sqn46bvrZEMC6ZA
oIttphBYcVq6+GzN47YvWtvOYAHg9cjTWFjQMcAJVjBSwsQRP0ZrcW6pN0hQK86ZucWAyXub8grX
QYxCU4t04UkYWsARrsDoESwZNSabWp5yfDxjWwTJPn6vVcEWSjQEcqLgisWeSnQZjnXAWLXOWtq0
P+0IkIfbNb/D2+4Jv+VMaBsdjQHd39tYn/cA8r6kwNt2OqnBGQET/Uw75tXmAc2mp0jvE7JZpQAk
QMm9ICAGZfpI83Lg9Uqkr43yXoNgqkGwP4RK+Mw0i0Ji+4W4MAIyDbjUnhThhFmmsgABRYRDRA/8
2ReyusmmrsV1sqLxKf94ebLOsGdAH6KNh2H7ouYcbfAVns7i3Q+mRA2Pe9LWdWytEx9cSxP7jMNs
e2oRc0yNfivdWmAui9GkZhJt4U/pDl6GVJzm1ReJvMi8kik78nwMkz4gNkN5qNEDwSjg8Ct6iJ5z
3LhL6lk544B2g1zRGLEdujiiGHO77LtwSMK/nTggHjU1pdwrZZoBQQl/1cxR8Ja2OlJhdgZ4GIbs
Y+t6UFLdRTtrN+179wjWNRNVWzOwjYeIXWIRhY9JD9Vlmozi+uCm3wCEmNSf9X3bAOLJ02UMZ5yb
y8Irp+R0ZBsIKQMEUYQOfKjlNgvDKorvlaAh1bWe3Pq05szMRGbHrlTSIwTwgblvfmI9xPDe+vr5
M0BghhS/yruNdQGuqUui1kr32O/bKcD3S5vOYnoonPUYdh6wMLYpN6GVa4dcc1V0/ZGh4Jm6ifXs
6qglaBo01e+wk5m2zpbRNimLNWfSzJAMp17uQxGJn0vJV6/b8reSpnBdhRvfmV2Ovw7L5tEy8Z3r
6OG0ynYlY+Gbpame7M1kfTJyLrKcvn6F8aga71mSvBWqyotUCchUtrOBhTAzzMtR3DdZl1PRCioU
2qzft2QbQ1IULyUyeHr11VgjYiZHaOKsJW2jCFoe0BTXy/Yprtfhu2OC8DE/jA2sMEQy34PF5M0/
oJAGun7ksPlspIfIEeJvReB50nWu8hH2zfyABxY8zcOuPg6AsqEx3Fsegs12mWC4iXDsCzEugOjl
tgMEEPcryEgzTMU9KVRf+5nT1fjhvRA6GJ2WsFfn3lKXNJXuVAWqvmPJvYhpBd5uhy5GT9psOMXc
OTyoeoMxli93H1cUdV2U2d4X/4fN4uvT8ElVpLOg7vkDcTYWpJoD8zChJhgFMhUCS7L9I4iZhwNe
5E9Khaa6728Pm0X+9QMN3EWKSmEW9qYXOxEAEepvhtleN9s6L5s4br13cSQcvz1loY7sW75fxeaf
1URwxEyMo9dmtOGcTaPvoQisSSIaSIgPGPpGVMm0Ddxxa7N8Fji09jO5bT2T3owyy4mfTaA9Fflx
JFgu2WMwnilri9G+gaPInq716fT28RocTiDA+OeGe7nthKimWjM8OtUNij0Ksk+5eogbZVIPFFOB
V3k5Cu4uhCWKcUzVVwRaUrSmNqpoq2HLv7Kptui4lo+dDYtkiRlQvNqoePJpAQn0oKc00GYQ/wOk
PMUg6vOZwgKJ4B98CrtbBD63y8MChpjxsBq+WlaZtVTNzz460jY/oUnwOjWpshuCIjM279g5gB6Q
gldOH9TPuiDAeydowwVWU9x5xtRyRoQcY78qUJtpHvNVyZf6Zqfs5+6AGmURObV/8M129qo1MmDq
CV43Oyc8DYvGZfOxoz6b6xBRzc9kT3XkNamRfK52DPXelUVJcLobz+P/LIZBw2JmcHVkJXobwo49
JY+AwPgG+TZNObh07hOgrUrHLQ0U8KrCu0euhsGRnKDSkMX8gaUHf9vvv1UEEfhTYnaptfOIKuu8
06YZz/U9e4a//nP8IjKbY9wgslvWbUVOtMcV+GBIhNdCPFBPAXqxx6ekiswDwnHlmMTUnAuYVFlw
sTiXpKuBAWArZgxAv9+2lV263R5LFh7/IFu4w7iy7WdEX3s2Z2etXkeIkilIVSQgTOm0wA6M5B76
xfU0xcBZJy2BHRlxXhkbmfS3JyLjKnqYpKTcO//ftolDyg4us+tkTyeAp00KuCxgIgR/4oRzJXXl
Rz0FwMMXYieDYr04JyzgBCkzi8HhS4HO964nQ3zcnOCi7RzJiCEz8aAn4PvGZ6SeyJzx7wzl9QFP
Gujvn8aDoMmr1NdYBkGDSDwj4fJOwZNHxAmmEZvhyv53Jj1Rl/SKtBJVpnXUTZRQgktPXnSzpaAd
tJD6CzAqdqRCGDk/fjWPysGoNmKvErAAwA5H+PIgehdvoqBO+pfcHkVspz+AatgmvldR9ihppWt8
M9viMd2FYbz3Vkcztk1sKK6ifnvQMxuNRU64dICQcTt/e8L3bl1CEHTNY3YLZ6rMBioSJ0uSkAxb
wfs1lcBkEdjQDirH52XoUIK0weVlKaev/U6dDsL2fgG6e0Ri2YogAR5j0bi8pSLCEsMHLD4qlol0
imcIwuCmFgRnZ9Y/M49quEWsU54Ckbvye2w+ES5qT9gss6Vocj7IcqGEApNwwmU5nbbGEX9zz0rs
6k61G4/247wImUfog7/DZ+vOJIdZjZzcfMDV6u/iuWhLlvYOAM66nUcWO7Dp7n+QEqPIqCeZOohW
YjIT9kQAxNxWsnQZcFkM0hiHuTA8Sh2d1WRI+SOI57v8VsWTziu8YCkUDX+Nvx8nVvaurMtljwwD
QRAR81nNf50pehyRZD/sKlHmyb/dqGkynPO4Pn2GJIyT95Cc/QmGTjqgJinKK6AUo866/3umzvg5
prBMlyZmhdv5vpDw7fDo0iYYVTk3aj+BCTR4iwy5e/44eVGLLLXcHI7LZL58A1Ecamu/Kv/WOKWF
VwK4Za5YZyfElu6VZXMhUu23DgSH9pgAW3pRHqmSrPvux1/r1tQWAgKi+Q7A2SLnxJ4YDHYZ89Zb
jCYMV4x6+pe60JTaRynalGMgLDa8VBYmw2KqTSvrSgmvYQoFJdrHnmbqpbxnfQ4NfqJj/J4jewCc
Njh5ksJiOEc/32AUDfE4MiErxUiDXwXFCND8pTPx617uLPCVT4muE/YilZmJIKuDcz4glUsI8URM
1Y+dFNtK4CyLd2JKG7QiBmLnlKqLoFFnLj0+9hJNlxP9TmudFf1A9rg+S1wW3ogRMtUD5v5FUUO6
21jqNwP7DVTQJshsQHdlRJ3hsPfS7b6VvsG+yNVZNAAF759VsAxGKuaxpq/d6Tk5qk+I4tyZnBNt
IxFRsQkpHleW9K2Ls5Q2/1setH5OudnxvWVDdaag7M9+iMds1wYh9OmnN+Czuv/iAIIgTS/0TMX+
JDlx5kWkmRVDHEYMyQF4YCO2zDf4Vy14Zy1+ObGV8zG6ro33XwtyRKF0jscVMSgHFEcRCqVMD+XT
NMjSgojSy1p4Bkt58bD/fGN+ifwkMBYwd/Qy0CtuDWgviRxzgsLPrhnQH1GTPZKHkMVD/Opgs5p/
7NksNluOPH66iZ9a2nqB9syzdrqcs+pkQTPhbimmaAfpcqjXlJRy50wowRc2KU901n8Mkcx0UTDx
GJ4dW/8oYqtVW5X6ku15VfZNLAZJKVq+jnZjD6soENESAQX0nkXGM8iPbrs1eWOLA52JG81qcA+v
FiZ7GQXpN0sExP188//JmLkgEyzvpDz3zfqMI9hAL9H1epItNNGx/Yt3Vd9sip83XQk/npLU+inG
UJYc5LNZnrkBvPjIFOtQ66RRjqJ+dFqJ7ARMWDGQ4lbTRexlBGQoQHt6Qut0UIJhAvGew+KAaEgs
YBHe/58vjRjwLcnJ/l9ut7KodGNHwQHB+W5uGp+IHHe2AGJwkKr+eGXxcRdYdDkQD7pPcEnz/Xzw
wlW/Pj0wb//BG5wvxbqth0r0dHC7vJmGI8M8h5Lda58S52cTCateY5nd/yXfYtYr4bZQ3Preu9Fx
p7jmyAh6ldG/c0UMzr/BqWWHEOTrsiTQLUUL/f1slFCXPTlaSf2OI1SN44bwAIJihngskXUXhBMe
uyd09YwAKNj06glvsgQCdQHLa9P4+6eMFN3nkYYOwkc8uV+CBWDX3byxYfNRJ0qDeNKTFyzMaFGO
Mh1PJ7OBDYIfEM8hnzj/d/AopGguyYASzK7JiScUh8nBEhGKqtDg+L9PN6Qta8ZfwalzJnnVdMOT
QFJ9pYo8kV3jQJA5HJ4b/eiSeTUwGRrKoP7GGKoPSQR8/79BRekqHSKyzz59dnzobXCwarv8oezI
ZMM6kBvCpfheZWyGfC4pldBgFsjLV1Eqc7nenL9+w6M6AEtZ6iLth0V2HRWOLikU7x0rrePifNTe
cUUvpyc6OuRJfNWifdwfP6hSroifJ2tni/o7VJY6vyLETORZf/o3PRhBtYWjruE9TUyidjTh9FSl
Ve0dXgsksk1pW/1t3ickbKjksoqcZmjcnKjYbkmB5khiANZrCZWB7bQkpbbJxPGcpy26sZ36VQiC
fVp0N2+L4kgGPaOPJgunYSvLOyF0ZwlJEfLR0dkKokVWwRri2NUdRF/QBSTKT+8EtN6ADv0KaHmp
2TMhfho2/NqDRna+y2QFhyEoEvQerYSfIGbE2ZhLkJZwWdypBjDECloZJFgnI/tpXlXuDuLDcID0
2QfEtK+XyHQjW38hgVLxVHRn0gpEQ4iLUhjAU5qaS4ERzPq2G2DX4jZmovjQlDMREqTdmHkO4yAd
I/wA/QjQYr8EUo8qMEyjafP0jpNRlUWm1POZUglxVeKGx8WAHSjN3KHYClY/klBImT6yAUTEWrnZ
6n8l1KwoZkp0R8oNsmQhdImh4ihGYk5smegI6DdtcOS4bh7z+AHJJeObDgNt/zQm8RYgJoZVOqMF
Q9+lmA1vdiGMO6u31lK5o+K+xqJtLInoppRnRrJzH6SK3ha5M8Hp75huu8T8Mh0ptSjpD03WwRb2
7NtwSsQArWlCfqh1jlQs1jnMj8PfxlxW8W6vXKpkQ5jP3d5zVgwGENP3pDy9fANsKE7rcodvumQ7
9MJJZrWsb41kajSY9DSI7MSKq0UaHhRAiQRpBOHYrYe+UONFa2tgtVY6lv1ZS3sk8kSeen9M0108
JPhVNK1u7l6HK3t8rpDLUe5f6b4TDrkv/bx+kn2lHyL714rV57svFGjqJ66oS7Fb4BgK8VsedPUb
vAu7QSir4eCNrCejizdLOdkLpFSCp+l1hDMwJRSQGEHptDRXs1UEFSOJ7U7QSx8z2PXeLIzUqOCz
FxBUh7p7FLuC4QnIW41x0jfJlSOxWzFwSfLbhNZ6je2RW5BCCWRiigliFxg892WQ7v+6RnJ411Op
gqN4agu+05Q0cV24ODBe9tVhDVIaWcSTZMp1xY5LfnR0Jq3vwyMOFC3wy2cIQpcTrolYM2RfWqEk
48Qb+TKJF+qELlEtvyBNSx+FUgjELRP7p6KS4HeFSkNLA8nZeDQnvN+3O1hBIVadzsPbGZw/Zn8i
aG30dqlpD0btwyq5Ciylvt+aVWtjQQE65NtWEeBgccTRpc16dIVwSA9H70ld1oQk2UsZzPtpZS32
Bvo1qrVu1ha7SLVha/LddQv3o7wlZaCSOh9Hl3AyHOvkrMvxbburjJC8drQmVaPZ34c92pYHOn8m
G1birZYzJQV6STHZnI5R3NSFAVWv2WMiPAfWca2RkWsPUZeXI7CzNhZ+Ap8WiMHW9Bf7/85wT9mG
nflN5UoBCBfki59rLLAjXlNtz0eO7uCSkcDMopZpe3RIiUNd91/M4E/Pm7n62sPQaQ32qA2KngVM
VuNdjWUhC5VPbakujwjl9aUUI3rqQftC9p1n7bBa5w7me6lF4hUOYthvjwBx/unrx1jgi6QO9kRB
yrEMGFvVS4MLr5Gd8s8vk0Km6DkJcG9We1e3rOMXT/Fz1mPi5fwtAKm9kfLHbU87jMZVrZbWZdKf
yzjYfwWOea48/U6LVVUcjcJAj3W/8FzY7uASKhlNOV/p0F6llWL3Kn7Ktmqps1ppyk6Vp97WnM0t
psdyYeflxri5metUhMN2/9a3gUBdvmn7FYJKJQpgJGNdo2CAD6fajpsVC0jfpJ+gnWMJfBFI0oLW
BRrR28yYfxhj+xmeUw5ltBf1enLwT55aLRgq6nAsAL3PlGvKX8ys7YAzzhMS39+pbZehbTVBJGKR
7ix8bl2dNqih3sy4G86+ij/b7dH1PLfrlLFZtSLaBaNc+cQ+n+T9pcHpL2WAXmrsadJvpxK3drs2
teBKh+T8b7fUXk0BicfOoq7ZOaVy2npX4Ee8IgC76i1WxirKNsjTw/DmKiO9MqgH9H9ZEnlzvDaR
aF5nd8hbArQADjzofngK+33P/Gs67vyKkh6/O/ha3/2IFd0A4UkbeAKFOm89kjDArtYf3tAHzS2Y
kkPqFp2CyN3dfORqI3MHDk9kMBDTNHIe5eAx0PUX+6jjBWxHNXfY9UV5z5s8X45LCburaIM9QTV/
GPGYXyRkwr1Q7J5VaA6p4onBV+WUzYL2uFVmc4zFfhIJpfNbwRZVYbOPYN98XPP5I1QeiCmJ85gv
tCt5eiZXwLyngYnQ00oYPyI+axzPs6tgG4R+PYU9wRFHvTUPC+51w8meyoTCwK4alXnJVOuV+c0A
glmWEFDQAcwzoDqF+jgwKiym4Za0zuKquqKo3ftle9EKoYeFFSnVl1pKxZGIm5ZEExlJIUxN+Szf
byPPQhTMfO7Ns3stuUwhCkqUkxnrRm44b9Ks+5PQvZZBoITvHd/TEfQa4l1z6fBsYjNZughBZmCU
cniT6TVQt5779Hs2siXqfnMf6ertoODe8zbCS/Tvvqzh6vTxXjvIhPNJ7ZF/dwZrCItRigSk5g4D
OD8aAJ5nhtPj5dPxGJEgegbOsi44e0SZg/DiqJHnypQ9QJwKYqXaRJzGQhc04n7B1uIiQWVqotJL
Ri972Pw0HQ4f6pmQlni+vSWNQ1vJcIAIh4vNmayNI692ZURYeJ6TWWKA9VcgUI6CKHH72kemw8Fh
EXySZZcud8GCYMn/NexCwZdWi451aU/GEEtF/h270AmiQ/NMxhweoYhjXgn1vjTsN7kyZOCg4i0G
3TSr9hI8TW/XhPPzpms596RulVEqAgfaQ0/i/UffFW0va5Eq2hTk0Dai7Pt+A69dz/Iil3PyyMIs
3v4i73tM67WjmGwng+JBzrfKNkNQdZyUkDh13qTcFk5OuEHcxIp3RryR9apqcm2PvzLhGJ/do82o
VGNzrbJGs8mCAl0gddG2XyM94mExIL0dZu5UBheJZ6sHMleDbcGdzuS6EwzG4uoN+m6/QuSkcewo
ohb1SSLDfOoyib0ett+DFCHopAogbwWLbuYKoSfErOQvg1X1ppaZrf2WrdW0cYobkRXWEu/mNqNh
71Yk7ITqA07OWXyLLZ/kqyFNI/0HYEnB5KnPeOhrYpCGy4vIHUxvmmVoS4b+IX0tUmJhre5KzGoz
lNc3XWEuHZF9tdvKaPDJ0pRnXUN17Y6riHEvDfISnbaZ1zZ807RO8FviKr0q9lxFEkQ4Rkz4wD2E
y+pxB+axSS5+6rVGDncSGx9edpfOA5OGVet3o9WJnikUwbO3rswVdLM0QwJYPtJ5R3mInd60XdmP
1c/aTXQqmTAwLWna73Hvpi8vrU5Lp99IMi3dgGMVP82gnaDPnrmrj14qQncsfP0puLq9DKUaAwgF
2f/4aJkY3sRignWCPo4IJ9sPKUybRlZujbsZEJhCbU1aGtnddT4p+cPyI4QpI8Qu1RsLhdWNK3hg
XTvO0BPaDXPOu2/0BgaP7A5xWnURYAneUh8TaXwO9EQ/8Bfb+O3nGgN2fYsLpiOLpgrNoAfYpVIH
VB10R1KYk0ppYCd3Ld71BlQZJwtLvyYb/xlBn/+/6XevrWbtwVWVrk8wF7BEFnuEivO3s6X2YFWV
EjrKiX+iaHpThJaBdo3ONX3DD5qzapv09MkpBl61e+C3xwqDq9/1uryfxYx+M/JatB4eA16CHz+k
FvddcUDPg6sCgNdD1RaQ4zOYfS/UgLspNHmV1mpHJ+AOVAfwl4TMh91BtpBsP2iv0fk74g7eBkol
p9oETIF9w36B6JSI2s82bJ8rWHztLsGo7akH32piW78p8vqM9NW2KwheXtjM6L3CvSXsG/U7rOpe
1Ch6ecyJyItAq3IlbUEZkGgE5pOKsZqVGETyT0KquGGEDIo41m9ybGmMKTBF2nZvkpyzXIVWj/cE
nAnmFull7BSYZvyC54P6wWebAfUnIK8os5iwOs1+3g3ho0UIOntzUjCvWHI1C7DjryQ5eUMWijIR
AgfBu60RmmAvy7f/vLpqACo01tNcHurZClf+mIpQaNM5DBG8US9HUZnX0z7xrkojqh/q5SXgZ3XW
bSOexXx0pa6bASLbT3Hl45sY6rL8NZuEtey/fPbjaHYR2lbq3JO4mM2DjsWnK3+wN+xrJbL3B4Vf
zpIbTsLuC4OJCpfltj9gS//R4BoVzhdrVtaDxM97npN0DAPW/1/HxepHIx7XGrLEbAV0DFWSyzNA
ixBf1mWjdkYiqR9v1BMcdWuyg7VKVK6l7assaibEY7CPPxhHN2r+ShNQvd/C9ovjRHYj7NrSVHda
fwo4MXP8O3qPU95ALelCTRfVliVsoHCyr32wtbZrWL62N4vkqMIOaTeyc0FbZVKb7WIqsokDu9qv
4HNHghnFAl2VVdFeWs6w4o7nc8B/T/87GSdaJ0XgKXp1rAvcYZ5twmUZc+AYX99QVWWsKHAgr5zj
UH7ayYP8502UbQHp0RPYJAqli4YZemIUKm1Ay30Ivs3TRAxb/UJrcHcdn+I+zoeUYkkmHM9d2sjc
R7lpTgYGtO5nY2A6lNbYp7GAsc9UmoO+BH7O9wqMofaJC923wecaI0O6hDyvOskfCv4+TpOmMgr8
NjGwL+SFkHAkxVvTwjSWamMBckFVduhnTktKHWBzECdAEgt5Rs9Syr6apuHdAR8qNZdS2uLGYsbi
lXl5SWEgZj8lQWgbE7f7GqLsZW09SBxavFc/l3Xdf0uKcFFqacRczXBfeTueL8U+tQm6e+PQDuWa
H2Xy6kQyLXo1gF7EbYCFLTIJLwj+vO8UQzAyy4yinRCQ3s6lffLo8/LK5Ow1tL0Ws/cGQ3VuuEH0
nEZnxLmdkt3bEIYSIwFBc9KLvoEYQTtuHAb3NQkg3A/XB3b4+qhC7pMgBW8WQvimmUpVQulzxteY
d068l+1sSDma3ANNEVr+PsXzrAH9bVtXAOzMRKjIO7j3w3ILGCLiPOWYuoEhUbcDAsgoRDM6uxms
wbszZGX6ir+7IPKoDpjNpk3siPNspWQncZhS8TIp/Y9HSjAxHNrl9C+MZd6UbKrGylhodzDNCwe2
Lw1UyNqM+HTTZyIP81C4sA1l1cDA7RCgh/kn5EO5tlMKnM9HubSb50i7hmUaKQ89Yd4WHHq9DsKk
yuaF2WLnEQ7TradqBwHTe1jo8/tXWy/FrK6TwcQZS8CjwpPmTI8mGl1wsjdZKhtL4Az6Qo11QK1E
L+RWvsagdYIbJZTq6xVejb4FVkTra7m0TB4THUC2uCde18KnE8XVn1GulIop5jS1mtZpz3pWtmsq
7Cfh445ET/MQIldSqDYIpkbU9YGNtaV/QxPKkLHD8AgqIGFm6PDEtGyKwD4f99Eaeb9CIonSg5yS
wTDWLVMy9tVGu1NBLbyf+aYmbccjX+4nPlvI2Yt+VCvZWs5grZHjsdQRQPdj9OOyUQleFSVPkyUa
2d7RmpWEehcmHSFBEfU3WFUmIdA1bH/C7OY+bQcasPS0cK8l4jHowVPe1gjPIy/ZpoczOiZQDRNK
dTVhMLBLNgLJwEP20/IwggAMfPp3DVF45T923X0NhxF6MBNtg5BLbvgqclNGe/asUzU/xjdw2Yrx
5p2NmEjO7+UrQAcGXNaDbiLuqwHkkjz0P8F3/aAm+vMbZfifEFr7QUKny6O1Ks6q5qk/MHqfguv8
vfLYnEpM1WKdvBXUoZQCJ+OLy2OV7BJVYzRCAv46L2tAmNGSXF6SRZsCQLVRAtiN85gZMigN3YH1
AyBvadc6uzab0cS4Xr1is4Mx5mVqHsIBwuDC81VhPzg2Ai8KJZIc7YYYM3eOW2QKIt1ciWIvEwtO
toJpkztfDy4kuV5M95WNcUCrzdSn21ssAx4WaLd8PnPCrRK8Dlh8YUohEEjY85ja5Ble5j3/YyLN
J9txQNTlN1483bKZ54QO2MmkcWVCU9JHlhlsZu5mWGiJYvOL2pXaP0nYCQYkyiHyU7dp3sfVucnG
vdrPAgb7esMqYJmcUkZcx2llaV0ShYUKgBusbjJs7oaavZocjSNRy2vBOlvsARQz5HEcxOzr6emJ
gtqQSnGhxGDM8ak6UQ5oOncCncy7G8Q93xlvymLLZ+1Cp23yfVGrItvIkNz7YX41coM8fpApZOC3
hmOdKiSBOggd0dcY5DqoEHL2Aey3k9i/BLXoUo21xhG0STRy2ey7V7v+fa/MUT/bTDA/LsCOF92s
2u1NpDMeJsIykaeYhdtnT3AAwyFf/mckST6ian+yJhphd+i3RTNU3wTjDx2PJd3LMXY/qYzhivOT
sg3dOUWTJiK0/tq4fo+9+ZqRzgRTkZVFcFvC/9ZoYDR7oMS0oQP+zVK64G7gOo5IqNBQkn/PCLyy
8i1kG7eJ6qOUdrHLhyrERYxAkLVsKDJavqzbyiXtUeJzyHlr+91IEPY8ikGT6RoOT2R4sCmhyue7
2zmYeswVzPK5cAqTaCwzvjbdmFCCxiovx24dt2Qmd65IWSAG7L3h6/onD/nUxWG3f7Xs3FatWw8X
MoKOOFBYHZV6Xe2gH4meo8cLBEoz3RofcXn/EQUhUEPN1Y8GVzsMFtF/kbpuZPN3iPtxBvpTnV/9
OGbzPcr8XQ8yltOL7NoSf8enbJI9bLUlbb+3s6hgz3zvjW2KW3K1Y93b8pueKLTleEou51gHyjC+
idZRViHBRTsJLIuv0mjnWcGQHU9/rU533fD66Wsx9DS+lwMImQQRRzXVee3MpfbaI170m0lbpvDC
griQiYU9h6HenqBHc0PYqqw4j9ZQrKt7mmi/C7n4MTcDSVO/TWE+02NhtmXuT95AItpWbC4XbSJ+
xsTbrqskdGtHl3YsS7pQmLPxa3y+IoL2fJDeg2BfedP0CbOuoROdnzHZ/1nINCgIS82z5mtheh+m
Pvu2ECaB490rWmLZfdrZi7qg8CvuSFXp7oaxwS5douHv314JGSW82Us6llOxHC3E2qtKcSON/GjY
qydsd1Uec06kXsxn5LT/4jdJmHV/WHQ6RUqXODjrJzhU9Ie9/5ehkCqpXE2fZmODieDP0utpNXfx
65/6psE8az8hcw2ShAUC0vu3AQfsbuxlqMpo9xsKsD/Ge6faC6HMsiuuuPkrJowgaCYNER9cKaxq
mau/QD0cfYm/iwVULOaNcybfJ9Z96lmzD49vzRnzCA+fhgBAHeFKTvMYS5unYIxdBZllAXHyBhnZ
7XQzLRESC6elxEI3+dDiUFdRN9lsMEnaE1ji1i+9T8eZng/RuYobtqGaBrGSC8MMoen3bId97i37
5z/H5kHEz/AwAiTf5esCj8PATwvrbPjVAEQye9EaJhd6bgMoprpAHJgOxC44MXMXG9lJIejD5DJJ
jlYWvMJe9UAyxHjz/C8BiDR14SEv7KSZUmERiMsHU/zD3kyCOLBqI38p/dGreMgSHaEJzPhivYHk
KSCADumHwPGyR+0X9oAe8CpDYWZjKJ8IIkz01kj6F0uNtcZbECHDBAbIwuRoeHix/+2edKWT3aY7
9JV4HBpYkzSLCC5bbE4BOk3QLzyjCnIiFNv6bnYsf0kmFgRwpcCzI/D2KIUP0pvKvQJrP3FVUWPn
adTZ6cSqX+hJA0407ujIhFCdBcwkdbjqGGcpFAlhZ+18ZyLGVrsRuQUfOEjertBB5W61WDZa0j0k
KFgsGqKtgiFUAO6gb1Aj9KtdzEzWKAJEOzhUKerE56UTqLLafxpFl4TVF4qyxuWraAx09uMAhq60
Kb5a1otSq2HWzMweU+1s3OW5ws+Kkai02jUyYMBGOUtzSf8LGD78HKGTH+TvPVDCmmkd9xpmkRMR
pz5rAZahJe2GtYJ+FDRspTY1QenbvI8/0OZdTz54d9QxhlV/qqF2vhImVDGTNBrvCmeEBhNvkXKY
AeCAAr8L0b6M8JyLVQPeWtAwTGdd5tAPM6px4bRAWKmuDlILSUxXQwNJHto4SYvaHlf63FlTUYv5
4GwF6y4Na3XlOxpbfKCiEY97xRxSv8zOXGD0l/wCm0bmXP/VEMVg4F5Xb0s1lsR1FYdZz/75+Wmt
xnNtVRsux85G5JD5pniLnSvjB0FahFbjswFlzn9qurNRpMPgHdlH3Bf/buZNCiutCEyM3jArUbit
fGYygG5xepBJ5A59GRBVQeH2u5+alnks0e/xTc/XJmmrwabXC8C2quF2LTxZTAwc1w/opg33wuOR
FB3LZrUeXnq9rY1VW/NwjauMm30BpqZ/9jWR+SJuNuBwoU1IcwVrwsU0/5aBkHkzhE3SDcm1IvPP
/PSUtbKGotMBkwk7/ew1awkj+sY9PZzMosxTKpBvAOfnRLTokVNO39q4IJkhDju7wHeCqhoUV8hN
V7CmWp/c3uWApr3gYkbph575TDNSneBEPw0Lsc/vZnje9lVh08wVycijC/W0AnzyWCEGw4sCalus
LHXstYRE9hDX2FkU9huVfxhVKtcy7agqUAtyknHKDEWu3MoM5BU2ReAlhkvMMBdtrASrc4FZIxpx
FEWXtRHfDvCvjcgNNG2sLHn6DdkdEBBx9rInRUlKWNkDlKCPOWyaFLMyLurMV0NroWvOBahcyCkl
bzomHV+L/sW1XJcF+7hR5OwXLp1iHEG0vfe0gqagWjE0blhQp4IrTYWur33L0QBSPuY+LS+iO9Jp
mrvA8UCvTWtZkcP9TqZQAfNQ3jkTjPyI+iI0JPaSVqWJYhsORsTVo6R89MWGcjN711ln6W/rP67t
qgvNY4HS1tA9yduA/oEcfh+wDpHFJpdYbuWCOsQx3doDWUxgIYUYQ7DObk/W6dnHipntGLuQG5uq
LrQss/zDgx+1wUbsXxKwgDHdZiGK1MU7XKOHTjM7PAvbJ7QWHCEDKbyv2d9Iksd0dBeJaLRiIJow
78vKAyWz9wTvBlcRAuYC8U0Uchex7I21BFeyFP30M4xiCD9xgNCt1dFPnlXwFjGYSYcCBmnZpNxu
TbQe494UU65r2lA5hzbY5jh2jQ/KJ849nH1awaelpEpz+d/ptL/rjg05dDN1sTqR1Nn23LKfU6gJ
6HRIYvo0UxvQloMkjV+BPCx21Hy8nqWoxL5cYfxVeXhlcBjWZE6MIyDOY3NEp7k6tSvdY2bMQfio
5nXvW25wSvbsaw6i6Ke7cz8LoyIraX0b4XMdHPiEPIOZ4E6rFgHWIz8ItNDVcrXc3/0oSMiO6oKq
e2CpaXXQiGpyXxiAexmiKoaHBayyqNYu0om2TX7r3cmjQ0o5h4h4PO5c2odeuXKrBzdwOpQwa+Jy
Q1Yn2SP8eIR7e8xQzs3VBkzaMvjLgEDIR4SIDu0RoGBEupqJE8ioEGZnIgi1JiVzmfFsblODLvzg
s/CQV2NPz4FDlMY8yuiCwY1/VnXWD/lUJW2nqMLTPuu0KYwyNMlK94vNb0LlnOlOQgcCf/4BFOKG
IjQR9fCgM3ag9YWzl6Sstsaso9MrhGvfG/oZrFC0mrFMqKnMEahGSFfDQFK7UU6pPtLkPu5Em/lO
nhubKM3zLTGBbSLzRFf/ZjQO0rH1sp7PP9rk8VRAB7pyT2ENrqjAaJiY61k56jHTWw7j/6JYta2O
hVPVivEfCH9u6xN3bdwZRGjqbYbEwtT8pB9v5vmt/FrqKh7lB2XqSK/WOgWQV2aaGQYAIQlUFqbA
66q4XnV2HO1w9+d414VSULQTB0k7oDBpT/FHgsc+ax4Q35C8pG8hszjM3vO9T587G3NHFErRTSBy
YlTG0+nZV7ShDQEJ2X35Qq+a93ERfcUaiqOH+0g2b5nHE8dsGG9XEHuhixLnwD8WO01rqUNEtlX8
Cq4N8bZeiy+rsRXVxQa8ND72/8k/yjns4x+dBq3JrC6g51hL+ub9tCzFhxYtaIr4chYHxqe1rk2W
8Tnqm/IGA+Ukw0PNMmFbOTPrjexyw3Zgiwi6Ak/XC+dbn0bjyC0i64/+abxmAxoOoAKJVsFZsEOT
GVhtNBYQgJRn10n9KEsSgylXKAy6qZZyKV2XQs1tS8qgZ6DWKoDPGh5QOQC3dA3qkAYJNYgRNwNL
kp5HcX9c2uKw9+2VPlco1xk0SKDSxkVNRDIEIIIf4uSrux2HmTKdVtkKdUksiDhurO5uHllVdO2X
fp/ggCisPFUkW25AeSszvAnDo1a7OhrCgDUoYWelZNxFDcKV8xyHN1WddqpCxhlYCeVojeNfVnNs
LJRWeUy4obi0Fm9MbGy5oe9hfmATN0t4GqVphl5KshGjjmO7nf66ZbLXJ0EaynL35UtgNqeNRWgQ
wiuNVjPj4xl5A0ySnG+9NimRXS1kiKKj/9o3LXqRBwo7v+6ir3SdSxRrFtli6jIXwYZiOb486QnO
sIELu1Ozlf1rwNBqmZzvqDVSH5FGmhxXSlIfo+/+0b3F1H4veRZSZYvljInBX3ziupjNyasr1zEl
D/mbNtmyVOUDz/fKdf4Fam/iIRGwz6if+t7IHXqxtiZNZCQiycOwdD1HuDjiVQvThhGsxVljp6k0
nW8XTaTh/2BZuNipsSqtwuFntnXlad3/v+cHlMXXII3Tz+eX6dtDo4oAUOdyLJZDLvDr1wxYXERb
7HYhpgMwVUqTFqLlY7t02L8HIOM9S5H7mxyOiyIXNmFWu+vXOWGAjANAVndWq4VtiZ6gRbFYE6EV
uGuBayqAOX3ZnSRjH2Oawm0Dzk9IBjkGq6K6DJS+KKjpRwh9P3CUAQ/EKTneSiGX8CCoAxTqeyPU
t9kMxrU711rFJwxJn1epQkbXTe38e2Zi0d5qFIbgGamNxvKgBlrLdp2TGji1E7u3LJUpqbO21Fk3
WlmZsUGfI0IxyUuFimOoIQw3S8UyH9IegsZLepuMo/hC4+gOQr7cfHEW0qbDyqgO4MzyYt9dmgNk
ZbJF7QxXIRYDx1a5GFEY7v2p0e+DXStbr975fDdznP5kmZLZgPClzUdR+MXowxGRv5ynAXVI2h/C
nru8M8coHI9ZVpEvBYSxeAg2G4cR2N0/3rHLuBwzQFuaaT/JMUvBRgBlQFuhf9e04gxgiU3KWLVu
Wg++0Z0sxHZzUwQt2n6ow9w8QVP1XKjryGXpqugzx3O+cGp36/r9q9AMax4h4/F4sqrIUdavB3Ee
bZEY8vkGUYDL1lrRF0Xe0AD1jE/yHjioe02TSKS0/1x7c+KiD1oFac9jA0RbzeHIaqD+7y3tBkrO
E9ilwRsQvYaP4AJCWoyADI0/SKmb+OM1+vbsffYoGooEg7uvmb950kdQSMhmTsV/Q+s3v6Bvan9R
1Ye4Sr7X6h+zulzmYxhaplmW9mAd7Bjn2oRYqlrKMvqqVCskZWxxAxr2NFwRAxPlG2ICoO4qsgY2
WXgqpjHHcTbFose0ry6ThAepbhVIjW7QVq974uaXW8+ZmHTrl6SPmGUz1r2M3TvNzzDiDpzOPDhw
P1TKHCI3GPiPiipAqKKsBUJG2HGN50CDgJeKfM+4K3Yxl88YGFSPs9ryUOqNTTlDraEp5Mo5GE7E
7qCZ3oLiyaR6NOsMPrQceN+HkEZp4YnLoFaFwSKWYionpJjXGz3YvOFnT1jdzCm/9dmgE0/tEx2D
zTrF8yn7wKXqJvkU/HYKZ4OcQYNSxjk5ZMQ3utLBEfaf1Q2QMHVeixWGrRDxbQlF9hjeGktsALJ1
2e9ogIY8XPvhlKceo4IYZoCkVHCUHBx2apBNLnx9KKAN5s6MAX0huE271AQ+/6RH40t5ISrzc+J0
Xxq4iWVptxHAQq0JvfnuXemCnelzwgXBvnve8iC9YvaBAmzcXrcvwLTqsgGUic9cRJ7UawbyiNrR
XHeNelEZ5uknal/NJfEeBFr0n/m4UmpbD43sVkFxFMb+RifnibhDicitLl8X4tiTnO7RfADrg/dJ
Fc5e8lebGH/OPRqFst5FILWeJbH/yUv+RdH7pfihHfoeCrCMBuKH4Jlxy1TIqQrQQAe+WbmoH+6k
GuVQLKZU+apOzlGcXy6nsz4U4r4cNwe0gf5KbxXllwsIjI+rr3FzGL0B040P4DN/IRsEGM6MipbN
bw4ADfjXoFE7UWi/7xmMnExkF3voSER/NyVE5JzRPD25omuxV5virWPC3rOK5s81wj/pxXT4yyuC
JAu3j1MD1xwMY1Vn05IGi28Nl+dtzq/sHaHq40O7oUKRj8nW8j0jjrweVj1LQn/M4gdFXqn0NNXf
1g9DpYtfgVLDLh/aRZGeQeYgrY7d1oDe3mfQQsiUAKEi7jSTRXbQct5rzEobA0bolZ+SA0v5BkSg
OdsmCGiVexxu+1ioM6peU0q35+4IiBfr6DCKB+8vn/ezHUynZNDcEIORc0CZ77GNZfsK5oNjUJ+A
+uG3Tf8Lw1xm8R7Sd158DH0s+tRw6nVsP+BkbI/kAgtU+PxcyDSkij8TeLkReMQHRC142JD9n6Fs
zy5h5vNySQdXsRsCCPyCX5i0p54uedGjQUqM8u0z8vF+GunZ0KPD06L7WcIfnCgu+xg7N7YDT4VQ
Dj96ezYxIXikgZ4RRASrFAtRjnB4ROv4XM+UIl8ZjsfSU/wfsyhjOzifkiFpaE9DXm53S3KRV4li
NDsT6EYv30j9xTNqHYWJRd09x5r9TIPDioIbxlLTcSgeP6H4u1NTWAb3FMe9srpuqakgvbLayQqg
nsherAE8LWUkkbnLRFYJRakatFAoolvYgY1sgbCAQzEcXTHl3qwSdBQTTBnuCDOS+1ByGpJEoDkM
3SvaeHz8e+MxY8kgZ9crrpzcw2H+8pJTeQ54oL2nuCpVdfbaduvsvGH3ezz5a9oudkYttNITnqUS
7bfTNs891DbEKcXzR2qLcmpPaic/redxXgy/bgyyd+cTL0eZaRWyTPty12W4avoNlfIcgMqRmUP4
WzVx2mKQdG/PVYV8QmZnnJuIi1nzydyxXAccE99OPi9U8YZuJU/meSZB/cC+dkVpmaKgBEVVyFJZ
C6ZaKecn1ijKBo17eaTRD2qLUp1Xmr8Qors1S9WbQ6CR2hCnVlDR84t5arRJsCCjRiSE5zZhnWMz
zZfx2I5terGXuPcn2UwkY6+29CQ1r2c+E1to9Y2oVALk5VSKOfa9Fcnh4+rn3nib4NBpA75TDsgK
4rVL8YDGEv300C6gKc8bCvjTR1FfxccaBXc29q0hED6i8aHFyWmI0u6BZDHLKv3hVZKK9bO8DO9w
+cPCizf2ZuEHzMs7NxQhDP9/ZaMPkSB9FWqOZydZ5MnzpJt09XNvRqjDc1FBv+c3jo/c6sQ7fNOg
7f/TJjT4s3oIximMAu8rJfSeR22Wf4hSmRtooMOIMuhjfcIAcIGthV/Q2LvLoCEf/GzZB0g2doaH
wvJJU/P8arOlK5REhhvrYn58exjyAAKyMCycMiydNNzThPtsgEhFuYIf3rriroAZ/pNnXdZghFAg
wSxkNn2Uhg6HwCudZFuwLpIHRL3EioKF2FTP+DDYm6O5vZk3FS/kJfqBDFGus0t//CX+j3QvdgEs
a/igb7LX0mUuYk28sgRdKln5cjWzkWFqPr3KXXQ5yjiHkLSBYSvzwdS/zXLd9mmLrhvyjZ3uYL4Y
aJvhn3Dr0sstvTaJqqdMHNCsiegOPkIHwhLACrLqUaxi1lzXBumKi0px2WQN40JshVszDCgY1fLU
GDOnJ6CBXCF/hxrj+j4boHBzKyQ9cRB2BqOyCT6tTY7Wqv2Itd3n78yOFJO3Vy/d2To9gbKyccsD
+Y4GVADta26AFtdQ60s310q+yL15DMsOFKQtCJRoQUQBsbgTlLKa/E7yrg4bPAoB3ujUbaQ0R2Eq
VM7c0LDH5SaXpwtDEBPLD0a5Cz+OzIGOGhVdouZisBTX8Entdm6NXEL5OAcKt3Ei1HrclsYgTRgr
ogDcl+g27Wzf7sPKL2GRjxIQn7lWljfky7PfhGyav5FqWgDbR0BPl3SqXkpLag3QQyV2ETPFCLME
/2Rwlo+9xzkqhwW2mzn8BcLwt0WYwAM8PJ9fqm5KhSXUeAyXOMlDkKVEiTmFJD2VJHQ8zPp8FUlF
CHnJbBL+b1yWpnrj03fUQ5U2y4jkGSEbIK1nBJ7myeDohvxdvbHKKTa1nt3DTcRJABoT5iEYTlzb
QUcxJPRlHGoFXY9Rufbfpi09bS+5dtd0I/41/eWe3ZL3Rk2pwhkEFmO1vJqNubSeMypt7Jcp1akO
UVRsCRr/S+Y4gdk0GUsZjDnDjK3mdPVNzFH33pi43fY02wSIC9hYfC8jLNHxChTSXQ9HIYbbITJV
Iy0ZYBRruasHgNJ/4bEmRwl8C2OuPs65TS6X7+Cv8hN4vq21S4178p4GDpAYMDraLX7PaWT8TZiS
8SV1uxD35xDfChGXkslExVZrEvd4r/jFA7E0nnSSe/4rAHZwoon5id310JlWdgzbxCSzzfqjIzH7
rmB2+B9I1tN4slWRXv/HX08A/OxJcDb17QYkdl5EVE4qQhjYniuVlH7cfAA3MK7tUTrMEIu46w5X
OWQRwPk8AVxtNe18Eooa4hb32K4yuAnlOAx/mTyKBNZRY6i0lMhu35TAiK2pXa2iNHr0BSFPkhaV
yNHvAMXDYMs3j1C4Lg437ifTQ9tXydshW50DEIIwQonmjkTILZ+qxnw1gNJ/mV8A+4/2t5JBReZm
TpIa9A3ljmbjC1/QpLyQiwHV6Ou/TbGFZfy5Qw0NC+CdFHXxoLKK94Nh/FbwGlG6XYlU5fj7stW6
erAuUhBFM85I7N3gozb4GaUXtdq5PE95qBZG2EXcHeODAPMvL132q5jHplhM96AtQ0NL4PP+i0ay
2GAE7+zGdg/YA5tJlHiHK6jm2anm8Rq00S6f6/JzSVyaRjqJ4NMZ+eWz8tDym3009+t2EawdIkZV
4V9d8vliulxIvue3F8oXHnxKcDzFr5ICE2Ui7SEixJoxRqn1D9L/bcYOKyYBLlBbgRABToyEuvcb
lTwBS+UhEEhm//Yd8e18+qVO2QvDLbZYcrkR+/nIjeiHWIIaRp1y51BFkyyAXCm82hZfC4ppifXO
Gk9ek37sPOwtKjsO7lKwck4WfeQgozWdua1MJlcwpvS3ysAQL+M3Q5UVRAdbTJ351dHoJp1obvHT
yuGfrTognYq9VYa/K5orLO/Uc+1kkq1Lzquim3tkBGka7iy6rb+R/dIFZvWJihZVW2MJEjgLa8Jg
8oGHLn0hnmqd+T8VhAnrHplJhn4T1SCM3e0QcpY09zH9U+njVQxqbTHJDxhpYyEicJKX7ma2lHRT
IlkOeYeNPwr1veWWbFJIGBzeu2ukNTro0EaVFjkZ7kqM51nhYDTF260lkhGYQYdQzZKu9zC0JqGl
ADRDE3nw9qg8XLztaQ8CwhccA4Ty/2etC1yv35FbWXzmECnwY9Xcl7oaK0sOyFDgXOuNzjmCYKpT
2M1mAclho/vg8t/ZBj6HRWQnMd8dOASZcDZ7AFxI21gXu7pfNyf+qv3dqc24tXlbwjEc1lRIu7i/
jadgL1Ldp669nLsK0Wjf74Y8+e51+SYtjXwobU/pwp3WRjb/7M4i49ZZ3Xb94/7daAyz9IdiQso/
w1cXgNcvh4U46p4MF+I6esbGtm73aY51jN59FynK/NphipuZ5ETrbIe0QBJK+IzCnwcwwdAfuuOn
jTr/HQJcZsZHqt85Znz7VqLROvlwP77DEpmYpfw2p25hMcBoGiOCkzQQrn7XjpOCibGrz0kjTac/
4r3xAFL3Z6ECiOBjohHmIdp7VLsVB9iEttjMNib8s5UghF3KTcWhmF1qMRGyA0Jxp5LxMG42mEN2
ZQQYLN7SqgsRYPGbbY/fgYls5SH8iIORkF33FiOSgadKK8l5l3zhYMjEZit1Bq4FuagdRiZ/OzcE
p0H5yGgBWDfVBz9m0RuajB8Mr4oiRt6HMZbrU8nMyobWPm1+WzZO1Luj3VAguLh6fe6wi3KlGWO/
ELLsHvvdL/UksIck68XQOjWZz4N3JkX8mkx7K3tmBMREqSEAXV4Rb/lHcJVtl0hXnG8QM8bDgVJ9
jf08aOgVlEgZhPxoRGsl0n65W7qk1v6OqWjyKd9icMx96J+BlhLwYI+mratCcQQTNrDRnTithvqI
Df5qYZzE2Ls2aGy7mnMHF3bHdXPFg1Q5ahrmdZ8JlRx5MzSnigMlV7CT8Fr1CWUlF4MIVtbSllMh
/kUzkhIPZe5G2L8LqMuwaYIVcpimS1YATAsLO1SBCjBs6FYDo6b5VEG+WYvTFEWzgwm9OtJTIfKW
kBRl0vt67VKhrcen/W43JSke7DIrx3WrNHGV0lyfh7m5rOPxI4CGl/nWOGh5RG/JpOwYCQffhvY6
RdrCVVzejOOlUuiFxBmpX64DN5OCYYNnG10AaVBDeHUKDxDTEc+NPhawbLspbkvM03TKJyVmGgwq
Oy8TfB/jQlQ3/ZpbHFk4RjoIR2cW0EFbsRyTSqcr6mWP5DbpUeAIJpNqfIm4eH+F+5h6j3Iag+ZI
/t78CfOumrB25bm/3NYC+X9Cz+UFW6HDig+424D3jTZEQ2016OR0BIF2xywru4q0xkbcXvRurzNb
NXLj2tl03CjxJvJbFuW9y32X8E3WY0dnGTWkGR07OmmlffAWax1jCpUdenm87LouSC0ACJmXjzr8
+2j/lMX2j+RT/UXmoT5N705KFjgGurLp8G6U+zTU6QiRzH0xa8YdJc7LnIEM5+u4KlnrMqLDymxe
Om08SatIMmIqas+1M9GoxdEGSCO/pA9Z6Dw8PHS9RaBv1sF3c7apNM0plp3FDMnPtQDmmHh0qikM
vOMfli9UeAZmd8//EP1GY3FpIewfaEN/o/rAMojAhkDspoPfGbjIemeGeadJsqvlLoTIW8uHlzgX
QVwaPI30TV3Ee//5nTlJNhB27m0BKFiYt/bntpCILSL4L2rIDosLxbTTcGLNLAUChoEaU/6c/GRD
laASOSiy/lQxohmmhT0pR580qDcVEb3nqAeDZKniTY6qrtwz3/ugFAlhPqf8bzyoV4+cQ83sSZtb
m+91ohYxzZSghyCY2Q30myOvV4s9jxU5X7aZ3/l94UzbDLl/OcQ+zdFFWcgd91Jif59eHownSB68
Aoe6YHhny1A0UO6gcKzpJOaTOFgepR3rsMe3lbGJUOec8ERgdwCClxh1ykXXLZKOIyoW8v45SVRI
Rc/Bt6SS6AB+yndakYNpv1+NWmQMUxuNVxQQ9+xCOgNRjseyhRZFyMXyKfLJQMcVe1xzrlMnaOPK
4/JORO+sO+IQA/maTHyWMGRzkFbgvW9nUgKreCW6Hu5XBvqQWefGdVca47Lz6Jz/P3xhqe5QeqMh
NG3Q5A73NxREkZKa+xjRulgro0T1nida1PvSDMmtlV1GqQeSu7drJjAAJaCGa1th8dPXH89hG14S
Duxo5iut+slieeimiTHmwBSrn0wTwUTHHTDeBJ0LmOXFjTSVpxdOMKlXFanwr8C8SG4GEBZAsM0X
BhHNj1q/EEaphrTzonyzxeNecKktpf44AQUYPLuUp8+VVKY4svDO65Jqjb8pSAsUFzoK9+A6dsGQ
KrU9qrhqe5z+VTtBxjQ/aNh+3HQD8q7OgGqjB5KapAJLdyEyljLc9KFmEx1Q25ZD9S2ubik9Y5+S
MWrOCRzNhwQ7cLNPkNZJ0V9tio8xpX4EnFeaIUaTQtM1o+I9tRy7QbYfo2VjIHFHhR7lGCiP+fxF
wPQaKebSRjqZvyMMfNmsV++bPOedJv6V844SXfHqxOfjoskt96B1GDuX9Mp6S+WuwLzZipyoVZtI
QTvQSY3c/4jDYlUlM5Uktc4+uJlWt7YjO2FGpMzjmEemoIRmh2WLVkMBAi56hVFI2OwgrNAkaVSL
ayT9ka1n6gXDPAAlMqqi9b1OvYIFPYjIPMi9MfnuePZ1PpbUnLZe3Gx2Ts7uwvFWR11alufeTXcx
lAoxWMvs7O5TAHvIAoTxVWtf+fEJJFA4jzId3QLpO6sDX4D3eWH6zfA7EUZz0Is7/2q0zp+gFJOZ
p+fdavRqAmhzFbLhuZOWoDYSW077e5IdKiUC9Mtq0M8xM02QXAtkMMFenXLU0RNXwG99NqxZnHsk
zxcfHI0rhIsX7hRGcg0S+3rzGMPb/sVYGRoPMGkvI0OG8JB2Df2RBnRBgUj6ewBycLAG88FqV/Sz
gQIIDV9ui1sQjQwoNu5JEt26buOOwUDOamVhzx5zMylpoO/da4bDsl+QXXN2C2QB1+rf1+qJf4wa
aWFR66X1PnlUVrBYq4INOxy9QD7yLqR+/sUQEk+i062W0yfwVcS7flXZuMDLtYIcGUZgTVrwJX9a
JUFt2VLZ0EdfUrKzbnKnncYC55MJyHYevmGxCglhEgnSr+OIS70puHTaTsQtqkvOfEofhEI/qyt4
zz3mRaC3vSM3RPgb79+1uehVzNxJ7g+nhylL+dxyw051lQW8RCJFS1kzTgRvO0G34t/wAJiAdgtn
v1P+zMV6AMEQkzdTQTBIvkhkjTFdNY928H7WtWKS2isShaVk4yuaKb8q0XwmwqWnlnMUr18N4Ohj
uO81rSc+lMx0LDZOsPyuGdsGmVd+5nZltIuZfeJ3CkpsOHGuQLWJYXHk9yvQTWm5cMvMyDbH70Di
qRchZ3lHrhlvv+dkIgPz9RjVcEKBtfOCnDpXHb3f6XNPLjtbHVA7i4wFq4dm7xX1J0rCuJu3AF4W
tiIDLDk/v55GIzegLcUaQgEUoQbHxlDIZFJBvNiu0gQaosY4FDmn50VQu6FtJoX4mf1DzzxZ+cHH
4RRpglYwgK1RpgaWZDZuRk1VwwcqJ9dZTy/Ky8Qd1EoJbLx5AfN0TZpn/cEb5kxkRU+TZqVscn6l
Chp1bD/YEZ59kTebDDI2x+610Xp3uBxLjpO7inKZcIo5bj1aRQl0OlsGvgiiJDMoq2RWw2EopbPP
MuPmdEsz+SqIoC+uAn2VIg/TqAu+oROaA94JwBTCha7xFfRMLh2ZnwnDpdFHozhGFxJnzBuK6VOt
Q9bq6Zw82BG6TfCuJuGrCz8hGTZQLvc7Rt7PZgd1EI8mTHFWzqOFVPnjMFcjs0jHStrsBjriI2sl
sJw/QEorTSAUErbc5nfv6K47qiLN4/HmfCFkiP4AuOUEyPtZSXvdTdHslNvW39APQJcrd/21zZsr
fAOtcg+BCoYRbRsn+ZSofVt78rgyY0+EU7x8786x8wcztpYnSTz3ciXACJ49coP+FNsUt6MCLzdh
1TQTm/BKqhIQrRijNATsgsJNbfLDZBgn4sjPiZwhfrAoU83c1ap1/qzhUkwFcs9hyWan1NNjj7kw
fx7tNHNk/c6sjb8r5iir7+AFmNu7JzJCrjM1Okbn85SkKaAavEBeD5rn2UmRCd4b4BGhL0Bf4IJ/
VwO1urwAaRjbK4lQRwJu9xd3cJSDxOR0f6FR7ZOnTaLOSAGXrxMXdVt0DgJb/qA7MzNEPTD5DKOR
mBC3Rfoz1mCPltmOQhxmj2H2BLalK8j5MLWdVcdUdKJn1EFRdCrQU0zjngqYKF38AaeeQssdyt9+
AO7mNyCc9USApHzHnPPC+/rqvb8vsCFlclisjA3DZCOh1V6DAioHmPH+gafuCyaqYcLD2n9YAshk
JvsEzqLMNlZ0wLGuB5C1Ls3zfa9HQvqPmTWt71vDWo+8jtSQMo/jCdO5eBCwyTIRYskP7Iqk4a0A
mv27SpfTvN9N6MidibXDAyGCZa4Z2fWZBJn+4Ib1lsMLqn1QT8zgWKVcFG0gzp7r2dqElMFZojaF
63b0bKytdZrYdbc6CP9rIO6MDPVrh0ogJhffjJBTfskkjHrjPPiL7NIZqGHeFLM8wPz4gmPnN3QS
Rt0y33gI9pdMb46ppHd44bcP99WBM1ZYqrXPSUf289GIDsy/QQIIuoXIirX136GJNSzjz6dlnNnZ
S7fZ89B6UDEAhdxOUYV2zb8crRaWrB3oqp9ICccZjiChM+ARj2Sa62GnWPgCc6L5NbJzUQZmad/+
Kkft1iXv924MaJlVhBQG3bk1lz8ldsOghYJ3hgYVX0Qt6c3yWgMTB9Nw+Pn3ZRKyBOZhmEz5I63+
Sw/EVNoOUdt1pN4d/QPQhdaEW2GsGc/y4rx4j2XqYMetsJWgvOq8alcgrE5f0OcapNuUjQs+1msX
gkHonMs7W34XGgS6gfQou9Xo64Puxi6lHlghT6DIQJ2y8OBrakzp+jTDR1vo25MaYyFTcHi7klTJ
Y7cdcXRVkp+6zYRBUMY+k0KPxJ3uiGGGH8V0vynDk6k9Oi70EHSJMuEKKy7lD6l3Da4giDy5n90E
z6365oNZFH9KRVVxdERloR3FbgEb/fI4NbdkEJkDL5ZV62J/0vHqT7VaTg8B/LP0Skdh9Y32sKr7
L3Z8ocdQEvod6tNRoYGPHnzoQT6TeiaRSD4J/myXTHkENh6TAuXBthZkejX+TkvXEhXU/eGRpYPa
Cw0WQYfKknEnZJSVH4yD0q7SBTRT3I40mgtAELlhpA5k4UFJ7NziT6UQjuzjuhvRhp+AQiEeFCGp
E/6trl8PZ8lADxplawk7nxN0V4kpd1meFuPIdMriE/JeU5Wx7VOc+FX0L9L9yk13vXlgTXaIQJS+
rSWNhNVPzfEiAz9/GcyOJVU3CuEHxDZF59doBoulFki31eHGpX03kTomPH10kfZ2zJbeyfbDtRBk
yPdIZeE0Dl1aTRd1ZQ7sWO+Akb3DhsbAhynUDJd9WPmTaPBCpGFS+pJ8H4O1IQ7/eP8cnGQHSX/u
wkcjSUyLwbmFhxfrheS8ip5OzFmT0Gc5ClM0XCovVwF0UQroBvyRcsLRGi4Rfm5eBb05ZvdOe7Cq
wSIEa1wPq9GXG02nBXV9h/pl94Hz9bkDwzikAD1BjwAoWbAUxa7YyloYiy4iXFhuzJRJRBl3VERq
JrvJYJwW3DwR8QMgSqbq7a/u+kt3IoeZHmSBS5+vmKrxfz7ue2auMNs7WKIFISpooTJ22mf0WUVa
5gnQAanX1dEkPAf7wwyIX2zdmykmV4IvcKjl03ARjE20fqP+1hpBmW8i+qZ8gDUuW2yRorJC4UYJ
zee2y1GtmuuqM4a/MJjA4dsO57/GeXgJmC1x+ckwLlLdxPi9j3Sm/w1E7vCy3b0i0o8Jv3lNnJHN
6OZyFgFSCL4cZZUNyH7n9RI0VLlknHIl85bWOGnZuryRnHyjg/480V5+fv/rguQDbMIOqzL6mTrE
2ngGwBHKIv8BUyufSwzjc0rmLmgkoyX7Rs/nRDoTolcF5LXLAqDLM+Rncf58ca2pISygFFzARTD5
ona/yw9xahu6JKDMWCFMTKSwsn4750AtZplrnbWSEER/nnF+Y3a5aXfbvRvseAjPzvYAip7EhN7G
eyOvEV1dVsyZjfz2t3NCFK/JoEwKbM8/zBalB29NF+YAKBXueOI25w8wEw03UAEWPEMtordGLSnL
S5stvVXe4nJOJAEQ8bJEPAyQG62xnYkGzVGlhDW1RmLfb9iLNO3jv5h04vWx9Zi5p5/lzBwY8A7k
cZEtGunYTCVNqh9qV7bxNX8itBj2Quy187u1aR0NNESYCWJUNV+uQM7lZwkgtM6aocxzTceSzPiA
i8dooDZhr60TEzK9z5az6OKl/ReWtTTLOa4aZE6SCLu9xLHqY+sXVN1tV41TRTersWTyemDroSoL
l40GnDxW1GBhqoHLPWAsID4zwBjVxte0PI9yHyJcegp+91i3sC45dyv+8T9U/7c8rk812bN0uhyM
B5uIFt+Vi+7c703FH3ahBz7KBXqon67VVrAm4L0HoR+rFuHXgO/Ub/LwjESblmYrNUS7GqYIsg/b
F4y6RfucI7AEcGxMu3IEmvem/gDqxo+ft+wrZUqXnc9/zkxCweWt4TMtgMRoVipYDzdy+1RG/5oz
kO6veqL1keBrsjFrN2/+rTe4JLg4QB4xBqqkI9i0ne53AGexWAJgg5e0Rt3VDosPWFaYlYFyE6HZ
/AhAD4XODngCFuFve3Qv7bdJCJiAWGNAZzpnzqJgM3HC+sLJaT4vej+Urcjpqj5ntTiq9DMatUf9
j96Ud4E4MDbKEzY3zG3aklhMRvMFTRxgH5s7wdbtE+zEnSrmFRcGgRYL53CztMtAPh2sIYmTDtkm
GWq8AITEn9ul2xKrCFt8IT8uJZHjKK48nV/J93v571KfyS4ukm5KgMML52jkOQRp+y24AmO6EuOu
ntsUkkZn33YAh+WfXxfal68yGRZ8mcuFKFsW6WKl/J9/CqzhMzysd74hAeSg6qukDg6s25wMPk47
86bwFpe16takKgA9RBX4rPjUJYzj57UcqY2VMauuN/h5HqM42Aak4VVLAlR2Ln+r1OTm2mqXYmjp
ZQzhI5sRaxqzxeP3db/E1x+jLfN9YRXsFKhxNz7GOtqnpfaDUi0sD50QJ7pP4JaibJpt9NE+vi8G
/nyp9lp89vYnH7L5Eo5bd7x1yckEpY2U6qgc0vg+fOFmcv4RP51dxLCNWKb11RaiIN7W5SfZof7t
YAKVP2PWvKb0tGdB0mOellO7DFys1mafJAdk1eqgqlGTIUEVAtkn7ClNebHxg3X14Wf9tAU3fA+J
2e1kjxFKhdbYhzjNJUfg0rqgGiEKA5RHivTjr47V20pP5ef3RFad4TCraEUK1XRL5mVvYXj2UoCy
2IjGeC/8eh6Y9JbiLc8cAFoc/1PkOzMM5CS4mpbLplvp1hVSGoSLnzP/xVZz6fwgScQuYtQVjdMf
ENj4Hu25JAUKVfmecky+Y4+dcQADIhCdSeFRcWvQKmD0G2fVwtRuUsRcqZEhJs94CyHiEys2o1mx
allhvcHAHrHGevQp2c25q3NioE6lDFs9UEEjZDq2XquAT9Tnxzp4HRgds2YRH09g4pLyLdUoSBy1
zOa79kamGmn+u21qFSsyu+R9naUyfuu951ah3WX1FT4ouejaZ7ASSk7FPcBnmPTKu5eianAt8D2z
lyvXqn5LQhZSHtiW43cLKaWozioJK5rMxxqXzNjPvhzBXsxtYbQ0qlfpOCFgIGYMLdIW/n6dssQs
3PLGFuy0PWCZsKdZOfx3FzMp539JIunPSq8dTF9iW0IvozfhPBfynqZ9hIrvxY/NxQi7E8PFaaRq
ziYRZadLb19I2aXMyhcLwa6jyJuG9u5trE4t2ivhAYE6C/EGaYA9TqV5jbyYqofUz/XdQql2OjHt
O9UqTgspkoSBeOpkr6PPH8Ll8plrgDoL+ZlPE+Xo9POWut/1Cn00SIC61ovCjpBvk+uiU6VCHSv6
/X9wiAzSYFvd5Zg/rCmJV6a/jA9pc2mxQhGqABtO9anzAf4R6fkw5Zw124ZNDsbcA2Qjlbu7l13e
jj8xDsgg1SAWlNV7KaKmiTGxAB5KXM+TUkhvi0xPr9Umwr6O+zr0RpvTk+jLUJfCNPGCIEPE0lN8
MH8umAzzcxiFz3/M3NgXq3PQVOvh7jqNG7yREnILesAVqfIofFHcBMF1dxWDu/LetIGxWWOEDb9u
+6l7Tw6N7HAlGNk08E3HYOczNbETthbNBIPvCcwrtLLBZ2IRqBaLoNDMjaUGbBcU6nCK5gMjF4yu
5kFMTg0YKtCCT014FD8xsVsXBjqDOWPIZh0igHcR9Tv3z2xXue5obZER5Btno8MBixvrC57D8RLZ
d+E3bs28FJQVvW6a7I8LUx3kJnE4KxmvTXIJJ/SXu48xo2WEPIH7YamPoFg4uAnslpST3y1haYiE
EmGZuNf8A/vT5a78JtcG8QshkbeTHa4FKoa3+xHnnezgI6dR21QCLQfw7Y6RUXC1QCGbOTbHgPCb
1E4U5BUigGok2rX4rBuCGOGi1Gt1Hbq8a+D0NhKpBpAcsLDLEE5WRHDnCzVf7x3lVQQ+NNGMRM1Z
JaH5pHIX4BEKRSb6UHjYUNVYNxU7dCwvfjA2mnCXNkTH9x6fKxkMSHASKD/SDtnLgIs7zmdQCcUs
XJ5d86dNkX8d5q2QGmt2gfzGGlOqvpSyPKwlkc2KKUzUlGwZTlU4nTQLCZMAzdMSUr+7O89MVlYr
aPuPzzM5P43w5aSpsEUycCG/H+sN646n0wvkUtqtWs7aj3nnRjMzvhdvixetHfg9ka5Aran0a23C
/go+hpoSvaTlosQqkyK9FofBTLoclEvS0j3woRatJo/+b1rxufgvw/X66UrMaxvu/IgD30LURT1S
4dBAOW/uC3ZNuuGRmnInDNSvFQk40/5nU8Gd25dEApHSxP8wWWVdL14IoziJWDKENaEUR1YTRnRy
+zca6vTRaxMr2b6z8njeNbmQYoejcPaRR+Z5+z3BG2qpJifRzb+YEEghbJv0NHh/Jbjctr4PWcZP
auzG4WwrIC5kFlQ6mtCL0xKTCiyEPxQsu+eQwSoCt/onxm7WUNOf029TBsCZv+ZwCMFcwxszmFA6
0o982JM+uyVSDyjoeh/RmDL63vSY0doaz1MjPEvCACCmX0XV1TAbzm2TknWCE+kZ6fPxjhk5Ltse
GdVZOx6XoRlRkfyc4rqqvfjqJ6K2kW8gYenO4LgJPrBG6YjfglYeYnMTlGoXwWLPUj6amwgMWI3X
hE4VpR1y+8At36oLM9AxweFSynZA2/jo+Gv31GNtC7aDwY/TBlbGkOl8M5STguu+31S7UMj5bFdh
j3cI+22Psrj3h+FUv61o5EQqiYd1VliAEGJDdJVXFnK/l1Cj6rutANmcNL9vvT8dTtjglv1FzCp/
mFHaE9aGv/xZAGgDbkR2rPZ7y47FSxf72l+j9/AvEHuxtg9h8u0AMuBgvq0uO30qpOd5Bozpkrhm
3cOMOK2onl5JHRzVhtOTVKM2E/ZKR4tlPlH9spdrN4XYsZOC8Ec2ytSZ2GFse0ID8k6o1/kbHiM7
kW27LYm81Fhr/Ox8R9VOmJdPm+cszTDPs9n+EwfC8gqZFlvNCmc+QslvUkBoUdRlWVV1Fb+JuMp3
+U9OY+WqSnFD1K2vsLfiW6xufezzyXJI/Mijpu+riM6nVj0SznCDX4kC9KpvsCoTnVSkMLfHbueo
3/5frEgm4Kaya36SQTLCH+gOcrnMK97xEskLJZfmk9IKcsL7qrFpZuMlWUmnHz3Hp53T4d8ahv4G
gV5gTfhiBkOciUuRU6Yp5S6pR3vmDgEUhAp3EXU6SsY4pxpsLtF+rMPWydyZB0C/wzCAgp1n7rrs
x8A7h/2L8z0/tv9cm2nyjFn5ZVRVhB1x6i5b1uZwLbi8SdyT0Xt1KNmZMCEbzHhyBWZaCIZVfoOG
VIIfs0Ah6uTIETKKKa776VkU4I3catAg/bJOhrfA3f9nI4XyTNlu/UeJ/Cn3BOpBAXMrceeK860v
5LPsaSOKQqpLRFxOpONn0Lhpjr8C/yoIxu+WwqiIcsnc8m8GBBW/zN2KRkv334lotoa8V20Mxbvi
tt0Sq4k0ykckB+c1UzOqEC0b3QOQLBhGfd8j4s9LGzBs7FB26K/bVlbsJYkbp3kaOz8L7VTIbJcJ
u3CcIblBMU+c/t+HafFCjaYm1sTpCosLsj48StPtlyPImxVw4EsGRmjj/BrNSDZqHjABXCgJr/v5
Wv5fqryvSCun4iwz31aUWdjLwrP4zLuZhSMf4jTgwR+jVwG1wekQ4HKAXVTvGAhmdGkJwMy+HJAl
oHTv8oHy5e9uoBDt1MqpFhb4NfXwkhFFJyKW1O+BL5JMRW2lTWGYUKGVrH3kXVA7Ze6dqfr1hs6H
eERWgjiEWs2ErTuUDmxbXcmTUhhiVA32vEdgDNiLCoRW6ZnItxfDPLcXO4247pjT9HqevBBzOvN4
2qwbAUAueYVvqPiHe8WGLouI3TRJNnaMU7nhuLXwee7+Nixz9fMAKNMXKhXOUePzBNqfpdiBAQh9
i1njctYRZ15K+WwS4vCtONtsEQFPZefdQxoWj/lTp4GA8zEcO8YU/K+AWqGvMWxeZ1VARQZYGBpN
cRVVzqTfLdE1ppsNVJ/ESVRzSkATSdTnptxY4JdqZUDuw/gxIP2lsbIvhEXUL9ylgJyI8MrDUAj1
D0vCTBsKHhs5OuqNnpWS6Lr1L3cNHzBOy1j9kN9ydkI/ZkRO5iWKothZRDGy1SbSKsniVICohIRH
dl5qq4ZxgigPWma1FSgW1pCBfnm8PKGBgGBmucG9MwLXr9yqHCcba8O0dOG46XvZuMNIrlXcdkZc
Wmq1WfUxlEoG1EpO45r9qfQIRiDbomm1WdmmKJ9Bm9kSmv2DTpAeMW+YlDwstXzvTQQAngr242kQ
a1G/6F4muePdhsn2zbUs1STeGouQ0TdAHBAWt9T1FesFzCUj0V7l1V8Pv8zX7aI/eJizFXo2K6hM
U6Fn+YhwlAORuajMyGmJahUpZnPXQsJeGt1oR8OgGvQHwBYE/W/XIc9HcnY1yZZTUy0QaFPneZXp
gVxbm5CPTzN4UF8PgpQNY9chV/M6d+fR+iSCVqERGVw20mic8yikrXKFkHREj0UFpxMrTFfAKzBD
7sf1epBWtl+Teskcss7Yp13vMI4YL+BOY/HE8sh9vKnHq/LE7eZnFmGtBjuVYuitQ4mgWEr+8pdE
QUiA7ZnLOA4B8vVIWlqMDr6y3nw+WycXKQ4hnXzvKMTVROoNIMMcVYiO8lZIQewVAvwU2Fg4hXAG
PPcacV/PfuA236r8DVHwdTTA8zQFR7Ml2tcvz6MBET6ypFVSDd6zq3b01Qvsk8tGG8lS6zBOtY+Y
utBtxn+LYfXvq3vTNQGBvQVXK4TiYxxb1WojRpJR53CU0L02k5xzDWea6ATWCW9vPUzP2An6CQNz
kG+D8Rk2mOBTmykNglFwOepN5SHiqXd+RGybW4Qp0ItOschwkptDNsmO/2tK1jJNZ6fO/+Yf0I+3
FxYdV8FHjcTyXfYgJ0J9GJ4mXwXU3jMUj+cAq4MVuAzLNktSHjpcMzjB5EXI7vFXJYpy/ScKGmLb
UKN+AYm7gZnq/EfR8nozRPeXIZxTi6vcK7ECbCswXjDPqylJN0/Zl+fQMyG3ISHO0fv0op4mN9B8
l9ZKgKrpHpUZ4pEtP/POpI9lAQAi7JOAN0pw9afT4vfU86T19hO++sxXAHrQyybHxrYVrtyCVVFU
4A4cfOL1pKeZN1Qs/V5/wAG2Xd+yDPiKTwxhw4TczCyL5GGMuqbLAsuW4TX3VBmb84u+g+ffMQwe
NRcmPHuFM21O9JZBhQhjggEhgkfwguC0AsXY6kUQHQtK8qT/Zn0+lyG+jlYxGYFihY9beH/22Ayv
it6EQ6kF2vWCv7bnya1Xk7CMvk/6k/BeTjw8QExQ3mwftljjnx7EjeR/GhhcnoGX5seXxKbbKtb5
o0rMvAaMDYQuoEg2b2VEBtgjGcVJLEtU33NNO5WEMzybZMxRGd/Z1PJ6+US4EBTCS5FhiwcHa78x
KmtvvmsLqG+PscaqP1AY6VfhKZraEoz974gOGBaN6tkRNwOQ08FbcR48KrcR6MzyeLhKbhgj9tGl
nXZaIrMot2detRSFl77rmTQjCo4X9x/Os7uv5i4zTsKVbWJ12tT5FvE/mCA9AzdYyyhWRZPlWqh0
eAoIeM16ZSM8CpwLFKpLUkouIKWWoq4CzhxbymABT5nlNgaZYrinQUU5JtYe9yY1bPqTVYyKMcQ3
hi4fR0lGqhIYq7cYx6QB4JWYad6+87AReqLWCwMVJZAOlDYvQ9pm2jGVVvkf93brGKTP2+OmoIsN
FG+Oyupiv1Trtn+2AqwJr2KoUQwZrB5vpyvJ17x4nGeJxR1x3GaIbd7jOSnzqEWkf+dWKnfF4ghz
zzE2ntSyoeHiL/SO+GJ3xufrzwjRf2SJGYN/JSqLfSN3c5k5+qsB5W0TRxVRHBpMFOz3wE/kq0Mv
bnZfWYlm+zHFQiSCimYoIMjzgSq4Dx3UNeP70aXpylU7swVUUTyfv0lQbB0Lxw8sefDGDDvaFi+n
0JuBF8Au6IwflofMiynLSw5+epfol1On101WTrjzjh/6MO/cjO0+LDf8p79W3z6k5VVUTtD2YAVp
5QQbMgS0tatsEOnSo0DP/c2rxwfPiL/SoK6OdsWlKElJjtY0ZDf5hd85MRIzWoW6J4lxqmlLqgtO
B8rGRXGwSWByRYE4Ku9Qu91y6m7v/lEplnXRNY1qmI7wW5zZ+ZtwfCm5ZML5diYclq2tyRpreKoo
0k9c2N4U7bIkDwV9OJNaBkM+ShEuC31mmF4tegQfCZIk0veS/f99KUTPWH/1AWw0uHI94JFaRPHm
yj09zJ0+gCnRsx5mr2GDnvXBnpIROiKjwCJu5qVgNObNh7fF2sZYaKQL65COG20/ZNikhawOwhMO
YdYDXQhS0JfcFbNhnLC6jOpqSAgAhg/UxNtzmXY0goI6gje8ZtpAKQDS2cVLFGp2nq1OEGk0Z7f1
ADQNL18T20zqTCS2zmDxulAiLEBFQsN/7XRVeGfzyXEiS+9RoQM0G+3ENMtQHCWuf45r2EkPYyNg
TY3xDCq5zmO+OBdhOvLTIAIrD33Ztu2rNz8GImCxt48DhiNB/UyxnkCPv69jYn95UoF1kWniqdtH
bwfS3wyL0SoQpZpRMAMoUA5vZe4l/HxFpHbqOc78uq1qka2ll3+Ns8yyzL/nuLaJvjSEnWoDOmhA
ffzhUGPBym5RQyagLsJP3jj7IbJy8pshAYiiKUw2Mtpwj78FPK0dtfAxf+zIN+6kpKaiizKPnBi+
wh5UmDpiVBeIjEsnBb/CUqmWb9QfGqIEe6lfVaOB608R8mZoQJpu4fSoT2ibaP2GRBqN6HHbPIz5
ObFozrTn4zFATYm12tD3TYeRCGlvCmj+foLa64B6fWcVEDyIayCENbAmBWZCdjApC6awDcDbDS4B
Mi3L65yXc8YJybNb1Apg7xtGzezgFSS7a6ecsZEf73HbgB5RcREaWPITNrMHiM0e3sWOR7REgF3F
6ddx/yplnblklSpaqXsUzZFPyXPKtBMQAEeX0Drpd0z3ec2BJ9AIEBMYmrDGubao/KA4umc9aFS1
AT2QXi/mLroDnzcqGzkcF8u0C0pIob/hC063hmtY/Ysb2CyEd76XOtXvRRmRCuJgBaja/TXIkecG
sE/v7btEbGf1A6+U7DUhmpmDRT57e4FJETg0dzzrJEJ1zsYnK/QclpT+LGXmbM64gizGOpvPu8Cy
LLFVD72dPwKayd3B9jU367fLAlG/2OJ2hU7XluO9fFsizqQ6qxnLsJjLhzVBdDwu/ZypyG3a2ZrM
Lin8vpFfdCnI9gsL8izXvxIzstYhjyasxTV+/5m+G2xukV/adM+HlrQlIDMPu1BWpqsgviTUtT/0
euIB6aHPBNPh+Lnoid9X0NPX2nbsN6OEoctPTP8u4IhmEx97YPbGU88ibTSmuiY2dLJR3QVcJ5z9
U3eZMBbHFoKNIQRQN3+5YTN27Y4s8qoySnXvl5GTa0eLFx/EsyzKou0ad6KcTN/JCNGjBnFU+o3R
cOYjAaLrgL6JlcluJWH7izTgaQXlpnbDP6NyDwvBuWUXqsazF/wykk4mzmFzOLaPk5yabIANMsvj
X0R4TNCtjG02bsstd8ku6uKM3mfezCv+SBM7y1GuzAS+WpSija8kWsHkgrvsEnzsAvOmNXY+xoeW
RSkO0VxoXoG32FT27tJeNuM0AiD7Qgk98/BPwtO08v07GhcVK10cNPRC32UKsHnJtFZOauJVYQmh
foxyOobNhwGw7hWlg863kv5s5yAQaXCF14HNhKzX2DeCcsmoFZFekBlHZCYmKvb3MhQ4Hhf7q4LE
ZlKlaEDZaEytXJ3Z6/sD3tny2hLxBWPKj2+6rypUrOj4iv6P8Ulike3+d3jUwBX7FwGi0NOUwkd6
+KghYkdp1mL1iuOxnV/PUPIf4AEDMRTAFJRxoERt+mkQAH8lks+rdC8ptsu/LmuwTc95kZSIiurE
YAnXBanet/BAbsHly4ekikGf5Fv3kP0wgiGgJh9A5epPE8YndH6PDGHPFjdoYKoDdsQzXO1qs/gJ
cKfqgsGlv1tBBIsmt2/Gq1v09QGLTOEovivsu2Gm4NEmJGkdQ02RdvMUeUJzh20caGMqsD1bqE6Y
4i3fxVL+kWPJjteNlRaeXRPckSGcuH0MXKJEb6RjHY3CrlHlllNE0Dm3i8k3cOX2zC0BxHibXG87
MSs7uqsaUs0MsL4tRVQk+yYe5VzVZTu1H+8lUD4MtxW5sZ+5ty7CIOtrpHHHoKfRkMbaavZ1K8M7
oRHnROTH3eFmPyXazOg0JlBnXfHhMudbs+B2zz4PYS+uWhMqttLkXlkQehnUruyyX7iQRpq8J1NB
slQHxdBD4exVgAGzVEQ5h9+1PAmwd6fvfaMywfQrVU+J8I/INibcGLSUPnDOAjobFoi6UKqrbymD
oEeykV9+fkzxkiLBdPxu+b8znyW+H4Qn3dZCudldTNGMxux6v0nuY+55zPKWI1bkoGWB61HKj/5m
N9FJUT6pTt47DaahbI0zA/WxmS7KYopkknLyuJH4bA5UkGUfEn+SLq40Y1wQF41uopVTUb9alAcf
VBMlwz9pB7CvoG9R4t+r/n0bvImB7xc8JgeTBRIfkRq7lReQ81a+9frVRvUCp/VCTcXsSG2lbmEm
mQXVVsXlxPyXzb5g4pgH4o+jyjxJ5cxQcswOO1RYp5djVS4Trv9H8aVfYT5VJUwQeamHaTuRl7da
4l9gHd7D+U6eAlFeP9IgIvxt/cnBy5wMcVtDebp999H2ciwGg0uU78v+ji/pXycQElGSUDyS2tJm
V0sa2yZAfme9Xz7vskSlb4Z1/ne4dpw0Zb3OUL5UOfGtL/nbGXSwChJ7A85bTnZ+WqBAvUvrQleR
xuSSeJqmDAfwZ/0CpmXHH84xiuGLH0ZD2JSwHHQmNxKShtxH3Ac/PaEtT2iSPWDSH/N9I4ujHwdw
3ajruC+cAEkSQsk6BCzmtub8kVfkksFNBr7o2nrQr1KxhyKt6GswopG0rCR528IP8QljAsBgfxrr
rdYzsJ35ckiqS91c5UgjQ7OrtjHFJdC80dcKuV9HSpo0FUbpqZpcWg3VMgDXpx9X99c3IHm9CDZj
44r+XEVQzNZxL8uTaEUJ81NtNhK2halPFV7LfwXafkUAEYZ8EgGzapQHCukEtIkESUYW8k9yiAac
GD4u08uWNWgND0TKBlbQsZDphLAHClMcA75wjLwNjwxQFYSFqxXA2xxLQ85LP5StAAYCclD5iZ/A
1bCLfm3Cvdq7q/hJx3mYLIFU77gs2XldIcE/+u40RYpFi7emJ82Mj1pUq4yL2eNuwGEpP4hkXuIX
MOXQEB2MKpER1ySAE8Jr/muqme1UmZdoCi7r/+MZAyPGCZTdYevtdGqHDmCxlLshWr8VQ0L2EM+4
yzaGtmohUami9KEJFIsDfjjYc96cpVsmkZhf7ML8Dc4WTnslqjOVyfQRGWGYX6qbE9l4xGef/XXl
WjUO8npn45h0bppMh6TJ++mL7l2t2EosXLvMauh1ww7MHsHLZ9KhcNGIgXbq9d8c75NhLPCZhohu
zf98TxooUDSs3skANt0mRNp+2TxQxhnNEDhjCxRF+7fZ2Wc2ItkLnCy2uhARMWH3AAuYlSwMuNJ/
HC6kFXddxoz6qlFKyRpzb8MKmfUuG6uoIyppMXkdLk2nBfB/3msdDw6J929YjRlWNf7HaimcDKsd
VmsbEwMh+IGzhoIDqxgeGbFFFlB2rQetISQ9sQCo8j0HcuYfoU/yfFeL69teyhrIee1U03P/Kog2
2QFVfUi/FVwBWBNrJXNXUDI7j+jOaxyItiBlBU5Fvttxg1tTHbwFKJ1crMpMjrSYC1zYDUHf6tQ3
8N/jWoVyj8Gmirn9ItpiIQLce7oBbhqmupkAU4Pw24SFhHl8TuKIujWlW6tBUPojSxylMc9GFYWB
w/WnLf61vt+fGEbJxKNJyv3DkFfVlw9caHQcwfWle20Sz/uGnu5hEAKfIYdDS1WgTGOVUPSjpBCz
0bKrJ7DzU8naZS+Sthl+smt9PI89+Yp65CCrz4kv47z/6KbTMTngLO8vnV2JUoGAhwmOvwx4eL4n
yuWK8OCv53LNnOwlM2pBU1jfnkI9kVxjsDzvTrWp2ocfJvgdOp8jj+vGtB7/hyay/jC7NuyCAwAw
pEd4UvCL1PnxiQtnf3xEqWsb9gvSs8kk2Gko2s17OE+wpQ7Nt1EdgXsn2iz8556S7HcfFhpKI6RN
VlfIvRTyhGfYPnxGylQi/k5cVOWfW2ASUIzQsh0pyCOHSOXjqvWfnTpcoed3ic2YiEOKXXRZTvwI
Mr9nRH8FypwA49G8X66N8N/t2CX6Kwg74qlnzCgRepuVoNqRxYo5sCR5nbErjg1FyuEel0fj5N9N
cNgvdvgAWyViu22yJmIb90UJV9i4rkSQ5tAd+WPvULcTg0McUBlXHl00fH8XI48wb7+5aaMrq/0E
hs3b0I73INZrWcym3EmS7kj66YLP3e8AYi1CurDKsuEMMK0YcTdDWl7Nu8Uxhh0i0udcT305N91z
fnAfEo6qhiVnL6b6k52hB9XzQygsbEuq4wo96JScncJvf+p/TmpCp0vyK8RfNKjq6A5o+bes9txp
X3fckkAkMptpFoi/Ak0jFybbDToZHa1bagc3z10vAPeJRKusZDPwZhKVlz5IUijxRPt92rUetw3K
y52t41l2MJF4OkE6ZtoDTCwK6+ur8zslWE2S/bbA4wzQVNEb27liP/enUJvok9BzQrzpK0wLgyFe
2EgNfhT0PLVnZDYKxWtd63SaJX7VU/JIqoSO19TLYNwhGOtkWf82whN47b1UnBqu2eKOOPp/Dln6
RNyuY4Yux0fenowZkOBzTqIt6QLLVzphH2+ZB596bLjJK+v5sLyldgfX93FZGETmDLT5mWgncuFP
5uzTxx+nUVenL0mV+EMumQ8Ex38Kn7SONN1alhWsi3PDpI4p3STKbLrH1ge5PEiUe1Inv1r1RYYg
IdHTFT2S8Q2q1WgdjDVI9nQYR87EtOJgSKRhiBPoU130MZpcsekfKjoWFBFB7ct6FqRowSCgdyVV
jtc5oAuUAYBHKdAyc6jzgneSUOmfU6TDNxXHGMdO+jioTUJkuv/a1BeHxbEM6n75X6Hp8fAL8oha
pIDTjl8HwtzPrKbWaffMKmq3boln0YmudDHBtSgBqHijrwrSKp+6jyfOsKtuC+0/+gLaYq22t0eZ
C6MhJ58umk9w/Y8xo7f1blpq4VGrtTPL2o42aHwrDCX8NmZmEESyrm3sV1siYropu9aGrsPisJzA
mMCMgy+dijkKyt/TGdvJXd3ausktbw+GvGfbnRwR7off3cO+RZslzsU8hgHi7Fr7dFpkIadWgevo
lNqRYYGADGwvGCz6XgYR5uOC5UbER6RgvWykP6WWyDwQ6Bh1FOA8Yf6Fv4QD4eXQuvKW7GaV3VHc
MaA74zgtmlEPM6jitcqz+lOUnMIi2Sfixq1fMBPD7XK8lZZQ7/1nk6NCwWqTNxS3uSwZ3vUBywW7
X+ySd6VJzfyYnEwWecKGGR+jnv1Cskmt2TcECMUOwj9hK0PJ63SArQT4e6NsJHPVxOsZF1COlq3Z
nGNJkL4XisGpn/+2I48mNm+9AMExhR4x0VSvaAoHHZgcWCzz2xboC8WTt3bzey/UG0eu9HOSL20x
4/z6ATM1+ZmxfzXOEGUjEwthNnRXz7SPFYP2+ZHuPdjtUHqpSoff+gJwANTfLJM9E8cA6wUSJNyZ
N13egJ8J4TGI9VK4ZA1GvF4xSlx8XppJP8zDJqOobY5P01b94F2UZndKZ8KlOTpa4m7ZA8FSTbvT
VWp2cFj5TBSFgbQH0adCwW+l9kXidoifO42iA86lOWk7vRG4Reza8s9/nf4JS2lfgorX40kZdmwJ
QqqJzHPnhW53J1fw59BIYFOhVeghANaE879ezt31JbOd/dYoS4iRqSFtKwuw8tR26h4+pyCSan0H
4cd629xjOWiIypldqwyATk4HbJMz5XnI9o4NX/GzHmATz7nl+j8Zo2cdAo0qq+gTuVGw94tlDX44
qfwQNpnwjXoUrbnRaE8Oi+AJthIMJF+AxDXzxjADgCtCm1nncU+rs6YdctGEMoEDq4GiNxK1A+kv
WWcTeA2wFbDlphvxD6MsP3vHEsg9gSOjVbMUNhitLVCuawB0xWPTZijJGJmtCXXz+bBv8ysGmR4H
651Xw/qH2tK2V7XTl63fiiOP6QCCrgJQ+R1oJdPIxt7nOq6LJo9Hlo3SqR9y79JpMkNvrBxZzIXt
X5Jei+BgTTVF9IGI49kXycQEnNBkZtlBp6xbQrG24lMQQ06RCUICKhqjYECLBak1E63Ls4g/jSAM
oaVy3F4C3ulDEntvlp/Od56ugKIirRbvQScb9EIVEBObU4mAUnrAkytWS/gJg2L0VIRWMXJLwwG9
gzarSpw+MGfzZ1TphUWCROVLH9PlXd/a0m1sWvtSNz+/HkgFYl65vZ/ql2Fy14GUB5TcLoApkZAD
pLmF+WYL9125MPsj+kl5EnK38NB/nQg6QfriukqTkh5bKoMisyA3MK0eSgVNcf4/e1fvt4iT2scb
UJQhGgmMxXgMUSuaG5AOaFpjR1TRb2aWg5j9Fbo3QvPVqaHCoVWUNgcJoQ6kuqfKY7ZncIoHFXtl
P+PAIvtrFzLpFnaTwJm+b+5D//PY7N47GX4SRmpSWozj+W+OdBnfbf/4hLMeFBeIzSoLsOEbTQxp
+z6pmOBlLP0i3cMhWO1XtznU8rl9MmKaaZ9ZPOk+1CLfd1XWmdTJUQElqCO1FWEhRvtYIlwGhCIl
GSkaMnjmZUNFPiDMBD3xHAo+nvrKXulfoHtAJTfwmui3ENHURtsRQ4iHIu0E1mULA4pHo8FeHin7
YW/OuP1YmY78F4M4T7nkPcuQIipBbiGDJLTIno+rrP0Yte/5ZuyRRcgsCrKNhWNBf/tu1obHIbe7
b1cZ7oXaDuCHgzrABupMCQPdHO+0xXRF+ZXik9cOmT0pztN/yKAfsWPFCcCcVFzoiZoLbfPaZTA+
2CxI4cvBgolbtCKulPvfwdvcuNrjA0ZlN7+8Bv74xKuvebTnZ9MySeseU6q1J9HAxikGDbxvHeQE
3ttitB3qDO/++fVN/gchquC5faFX8E/HyW+Avoht/V1C9U09S/m65Xp3fmIHGlF2kOhxtr92c5RB
rfUMUgyz/NFtnjML1JvznCS7tyOZrREyFiwFpXCSEMDSlonaZd70XbnHrRv9G3StQHZy1NUK2HxF
O+BhOVl92GlzWvYCVj5i2oF6xMrFenG31yvthB5/RkS1QBboYKEhvT/HmzdVkzphPIJzEdgRigxN
Ec2gsTDr5IZobvhpEgOfnBxRQM+MW5UgrZqCSAMcPf8yUcL8dJF8VBd+hpOBXKiFXvwU4yCf6BOE
WSaZ5Ng6is/kfz5v6FxMXItGwodhsA85BpGoUkzj5cD8Jxa3V++7oohkV2lXP5hgSLj4Rqkv0qMr
hVp2KCKNiG8ojOo5rLFLG4sk+oMgA9qrs5eQPDTk+DicQjIut2t6HqwWky21E88FsFWeXa3QDk6h
1AZBiUsoF9WYNLaBwseOnVAxQ5l97T+jmIfIh06a7NCrdPpdYxMLnZG0FfsUTbDBXBebOQ0hSlaF
aIrpG6CQrZCMHkitKoo3YqNbA0oobMP3tpO90qpe/IR0HfYuBl+7hAWLSFCTwUAbjHpBPDZL2+gs
RylJAXdXDyMmfYr1Pi4/vsCiz/HFqqUvx0MOS56EWKGq5ps23vlZfHKUe65XBpFfIkJm4iKRPgTw
0uWdZNSQogXaIJ0MVmHS5iRuiFm1gNOrLSlTIFccQiJ7JdiEGKZdej7AjTaBAtZD8r8cblpLGsDj
vt4cabC6jmcyjhRKmsNFxbxMrjifMkg+L5Se7GD1mehuwfWZfISg0Gh1001zN5flDqyU7q15CIok
JU0/x+Ypsu5Va/qY5tjw1vruMDOol3F6yyqmUtiavYy6f43Svv3BGoNu9C5hj6dBL9Vd6GoOFdwe
SvJM7k5KZhTmjr3TUbLIljshOkgv8dlaxeZ40i3TQ13u9wbKCbd45Qh2es3PN1aWr0Qqn9wTUKOJ
ZXCT2Gg9wXT6eKyQx5e0XiJZUuIHMw5n969C/xfMc5ZAc3WFDipFDkbFYtd31lOq+LZar7zp8mNY
/1MMlMeT0ej4JBHrDGYrOSO+Z7NTgdDC4mFCswTXaTa9N0eHSZ6c1ypW8bsuYQ+F95OsGga/LxKe
e7UJXO0E0OhXDKGUCsS7SkWh0xNGWAnhLF4ah1QTkBmTLRB7YbzpNIzwxA50y6jAG0kmX74Lvtvi
EGG21Mw9G9hMLfhGzzKcu76T/hHRU2YTlgscHPI9O1hKicJf3O8X0fMrRYUtqxKfK04gTCT7nRgf
vAzNw0wyqbWSU5NS9hqGWJDXovaM1eL7fDty3xpems0bRqRuaUGzYdpBFunxLRyNB34zTHFzEeOP
WfovBQ3ejlHWEzH9vmtoeiI+xqYIOsvZdHWOtZTrS1iIwXZPnYTxOdCroZ7R4Yp4PjYSqU59MtUy
Rrog6CuexzdYgPndwFI/T78DmK26MJGpw1z7Skq9OWxcioTh1kh3MGlRmnZXWH59O0pXmours7nX
nB9kCRXqxFg6Vum3yTT+KQNMpCyc9gw6rv2Yq8Gc39h5rxqBvm1ybLn6KuL+Dpb1J9AoH9cEQ9Ni
82wYQemyAU6bf8jxDh1+2iuwmzBD+Co/VntKgMxngJjhF6aw4Lf59SDpRoO2NngW7HMYQdt46XAe
Wy5T/fi0W1qatWt12spxpLaEMGjG/G7Jse+x15iMRByAlMJ2S5MosjguGUog/r320cg+yLQC/r00
EXwsaBPDv0dXHZtDzfGhunkWIJLdy72QssbPw0aBQM/KMjZh2rvT45pTQQTtjtwx1vGJUbaEaf2g
9C70r23CNk1xb7agzqrIHnn2CD/0WyCucwvPt1LK/u5aBTMrKFsZWPJl5HIgxpeBkoOqClskRg9v
aXiQs0tO1Fy5XSmIhmf84HwZQX9Tye54g80XBCvPwWdNA54+b4UfACOWzFthTr1hJ/WzIG/Sdya3
1naiQqaOI5Lmun1d7di568nIr1uKFwK4tKhB9m0zHwo5YdLISMfSMmb37lJSfEgHNhjAT9NtHm2M
znnf/3kGv91Fo/fEC5bSTqQDa9zytgvu3Z1Wn4G6n2Vjnk8fqOB5r57WTl34GcWNKAXjPOfo+tlv
sW4RQ+j4ywmXNVRU1PI1zuVsdWvAtvUlwy4wxjYqMwSffW4yn4LW3mWW4Bd34bdIZJblactONvLi
4oLOM8MjaZ7j/N2nN9HXmSZRiUkUZ95K4fdNrV2DfjVbt6wNA/+x2E5hiW5RghtSxJqZyYVMK6/j
AsAIwg/eZr2KhMVnXUb/zL3Y1k51Kx8wai7HSFAVCsD3F7e8AQy60pgGfNldJDpfw8iMCoxfzJS/
tGyWJ2b+7P3HmdChwm13vxJAqnD72hcStD6gB1mi8ArXnSLuxaRTUQREkCtlIk+wxk9I+i2A8b2M
ZYVDUUn58QdAWOhISK8WgN7+ZZ3dYYTN6pqQhPTpT8Qgw2UQbcop8kEhZ/A22EgaJGxnyMvCVKTq
WIWbrWKY4+ke01x15aBW4nGcKU+79AxUH3J7AwK1Nof1o+a2ZfOtQ0KMjiIiqiPKS4CaO5FpHfhT
XXGdVGHf8tM+5/AxWirLtUwh4sLJ3twnsy/FP7Cy+eeSEkwsDm6WhCl0CEapZfB+sqHt9Tzurz+8
t3u7YfH3k+6ccdfxZ2r+Tm5mNbtp5qMe1wCvCYFuF1alVXnCjk0y5WiUOHJC363Uu0TF7jv5KuyI
1Vhcq3awjCtpOidz1vEnF6DDM8bDpswWyvZhUnMigInEnn1ms9dUNvh9qx8UAIG/O2X31TicCaWw
DFUpIkNXCCjCJZI4Yozuj5CIWw63d7dPppl5McZXlM9F/REMHnGhQk6Sse7HnQ3IR8OT3hCBH6VP
5YYHeF/Pyg6R9OmJnm1IotRPkjTDOlBeLD1Wymw9S5S0clz2e91fjcnLnPoSh3DhPq/ASs8d4O9m
uHD4PxEU05euL3U+W/jJm6D0pcpL9xes3TZhr5Em5VRZed7rgQZ8C2JgmcoD6+dmxX5bJIh85Qng
ZhEbsDuzDJ0KxPXrnmIDrfecdbKkSeg6TO3DLO2WN++89gJS7S65X6qAlSaBcsPtDEdqEwC31/ti
GKLbUtR8lR1GFxrkV3/ln47Ayynm9ESnFSvkQTKtZmfcXyqFSWik4huKHJ2zWaCM2HVuSgmUFOmh
U8IrXie4No61cs8Qhxx1ZcGDnT2xNrC+j29+59saGGIRj2A0boU3bQXznxIEY3yV7zrHT62FCn5b
MsPjXP7CfE2tNy39RiamP/M+yHOSLCU9aFDBHgV4USpjtzPF5hdTt5OCY78PL/Y6gs4SWCptqjq8
GfjRM5Yk593Z+4KB+U9+qoCBEz2yNhNpRZl3e67z9J/kAiSkgufbExGQfqaVLy68x+gX7c/QiEWI
d7imW8yF6Oaiyn/hVKyIDbWQ2l0tbDdumJ/epORH+hUfUK7rbh8OEAKZIiaiUOU4XG5c8Z+DlY+E
y38gXlKUIxVw/9MufD+/S4JJp6/UmrKl8eaK/mT/uPyDsly2qtSr0K1rirIEaiAqhze+HcYtxjlu
MGV6MpSTOqEKPuoiOgqRmXKcV+jFKrGY9kBUQrvAIwTKw4bap4Q/W6HDZdsQei2awtfjwec11CXP
+DRhVFP9dk6OEKHQzRRnCh+4BrqORdjheHdQgKHW+oLYLAN5M0X/v4ho5caSXqifGfVATZoBVsPr
X46qQEwZ8hc8+8mxda2ligcPduERrG6UiJcc8DMJqQwcE672/SNsAkhS50vC+ddcwfITf3kubsqm
FKgCKzRN4od6Z/TI33/OfEUk6z6+PXbQA1HhpCTuwmzjD0LiyTi12MhL6qiOh1XrXoZrawHCk1gx
1QsSwvxphbq1CP3hxLqEmtZdr95AW2GZTYICzmblX9P6oEI0DETLhm0ElnnOJmZWpJEukwLtVKv2
DxRkdXjGZodFz7KHV5GnW1nKHyuqfNG8yyX2a5CrVNid8kAaghR0IJIKUaqGkHEpeeO0O+CMACxx
KQokaCt/BNy/jnO/R+NsX5fdLPeiPSnBWyDO5YFrvd+wILbwBIjAIabgHTe7yW3sU9KaSnCldYAr
J7N8dtdZQE9i6EY+rddjrTGyckyGoX07MRcWyrPxNOEd8ylHoMcf+AJ1cJUvMO7Ut88Z1qeRhdRb
V6LVr24EtpZqkq3A1tM9GMp38iC0M+0FGMAE5ugXesgqvhLTskTWbogp1BooJrQOoPfxrYLzJw29
wgMyijlXyj0WmxFUJNafZLBrHSdnpqGv3S1sqH+G71lpXxKBTNBQA8B39dGlV/MHEjhNOXTAMKEH
w9F1JgIgr7+9Eqjp5tbCJi+UjSB+V22hs0Cj9eUddhmQt3CiDNzdKNRme63BW3dRHScYuAdoffh6
qoAm6VDJ0JQshC/++qIhWLxiFVJoFjAjgarqTaa9Q0TEYL7GJ2sD0EfFDYuenHFbp8PJcrxrpLPr
ALxMHrz7MzCH9oeiexfVwSvCsklIdy3fz9L700KZLNkEbzky+5JPjmwCBxOLNX1/hNjhZT1jbSsS
/v/Cgs8GThO1GLOTfTZNxUgjylr47KO/OgKs0ZsjJlOyVLq3wxXVZymUAqAsMK2DqaZfW6IOcRf+
JHieAjZznzikLb+PnwjdoMRVC27RpbjAVL7DNv040IAR0XgyXugJvb6ko2NQC7mnG97qeujJFYJx
sopRNMUUORHlS3XXAAJvPKF59AJCbDzWxxJt94UfKCjfGzWPyRluO/dTQbI58oyDmGh4BaYFzQcr
Sb7q30oTHRHpzZnNDaNox4dqwJ1frRePjA8CZT8xMen2MUgWDXiMFWYiJOEAyCTZnJL/gAf0/zbo
VUJK+cAke9UMCoJtXg+ky9dqpYbDf9+betVu6bDNhrG3KX1wb6tWWODGWJgfhdpcCFavfQqMMI80
N7tlLkXOjDPe0wP+MJGaazbNwuVXwcOvX1uZSV8OGwvcjZaf6iIuwqDkGTh+J9JZrXO8uaRPpS6P
too8gyW9XinfwVqwyCtD6/Wj3CVkhP/yi0+g0ifmZHzqXMR+6MHf5InZPlgxbk2tMYy7XHQKvMaY
0JQIOE5tiWvvKOq66YfcmM+oFlcqeOBdOgB1szykD1C8KEsIYRRNmnq+XLOkpjmmKJdJrnWOtF6y
sc/AXCUMR5IgVc5TGsTvMhlzy8uMGK40wBAucie6jxxLYUzWEk6J+skHNEnNaPYyEeZ7dhojZi3/
zcsLHWMCrg1bzR6dPb5hxmwjavWTqbiEXSmTThXctH+nlwxDKQxLwu0LG2K/lkjbJ1y/V2naGQY+
JZ/iSOgsf+hRyshoXVYnN1APrPw4c+dCuB1oWZBFwPXgR+9+OcZm1rYqNhtzBtecvWSTHRe+2T96
xnXRiiVz/t2AT6degftL+4tyJOtbRqgEG+pnc0ZlerGSPZP8YXyOyrhqce5kcYgwFxJ/1kmrDIAl
L7NlJryuSZ/GzNz+Q/QVbkSJcj3/dKwcy457p2A9YZT5PEgsoVZ1kpGnaekUMRcM8Mg3Cud9rS3k
fKj49dWEUpkUn7wW85HWvIAnIzlXLK5K00e8O2lOcG7e4BGEelZR83YkFUozp6VFsRx98H1FrhGL
wTxSBKtNC6/6Fg1q2MdfrITb7OIYA5rQz0g2rFOb4KyI1YMa1WrMKG7WDGViOdHkl3i0rgoTBtLT
h3U+TRLTwuc+34Fsd/aNf5BfcXcqq28gFKcFmy0QJKz18Wk4YqyJGR0TntSt2nYKwEtgKIB71WAe
e5NAY5soAoFSFSbWUk1kpordpZMcIbG+tnkeQYCZeAFqczRdz2h1up72dp3b6+/P2lWvdZiDJeRH
hQ6xzQeIKlxlUQIS7oMQbhvdIsJOPDuj1RbUHeyv7mwQGPPy24daHSpX3hJuO14f1hCTpXaHkLV0
VQ1LCK1S6lB9FMJj0Xfo/IbZTrXCrfzVSLcm987EkXlxfsSCf4ZpNeZelIN8YTdjAet45ciuyOse
aujiHcds/pbC/sfMVnJL/RUSJK3pse80oOw+diOrpP+vZDcMgApf9cMDLHJ5hWPPHJuvl7dEpYtb
WpZrVVJK3/pNrnujZUUNOJ4EOrNYHLaMflPHhCibIBaMsyEtcMBHmjXgCpm4dzoGFIZSj6N32YOg
wMZ6spVAsD3pjij1ptIyr66wposfCjJOaaI4ItWaUXh4ta+02fnZYXT2m2KJaR8YQUON7GAT8Tm2
JLpCebf1WADUOwbYWBWn0LDnUA6kTrE+mgEpjCs43CjKU/iVbp2TcGwlZPHA3m27TxSfIY9rFtbP
A0deJf+VkdSYCsxRp7QBxbbYAoC0L96MC8DJpR0HPqNI3nBs/Ztj8zoklL5/pN44EBvfeGq4Di6C
7kfsrqnmrYkML++RVlMEJd4iQcGZ6mw6qWgqcNoE4ykfwRTmceIHzqmY9LiHZ1mQy3dE+zjY0Th/
T7Zby9djhqzxV1cjaIP29gVeXzn1Y2QmQxyscj9rxOP0LsySP2LFNsHOGPQgOi2fG6U/1t4Lq0GL
wzMdFd0FREdscKEWTwIg07uH1ygdsdMzLiUMY55wr4XFgAoY6GWqZZkGzF+SVRNiCBupSWJ4jp90
UfuqEwpJqD18C9A7staq73KT0h6dBAZx5zZeR5c48klv5AMIB+wabpvG/oNivRXOaW6XPM2XJnTw
341jlEje95w6t5TRgwzfKFzetWDqvwOi7J6/+nScIzC1/O33uLfvi6PA6kwLtyVk1gF3HAAxt7vr
q0WY5doJZgl35NsExUyx8O5XnXfOWW2fnuPO57BPjcu2PGJqMljdyYZnhW+oiaQ16mtKPzy+OO15
UCkpCn8J0VSxDuaDfK/H/TlIsQ3WS79f08cRTYUIJtMavfLlNI41BtzgmS0qu55Mo7hV9SCkwV0H
c1K5NoLJhpxNBr7R2G3VY9gJaxGgnjPjbpWjygC6ofkPbIZcvZYwB0ZXXcl4T4mBK7RRflnJHVhU
TPenDcPCFyzCouhB8cvRrN2PtYbTKnjrITPzCT8kHtgI2AGBSb+/IjW74ZmeO6jgDWOjeyWdD5ml
ml7wh9gSmvMPgoJpdgkcHzUdzzELtmq0LXfzcfQKlLXs2ED3SIoHkUE2XUBMpTXPClCERzpQgUdA
iqzaEZOb9z8tiO6UOqJ7XLV21f8I3BDpZ4ElhxK18eRDAaAGE9dglThJor6zOeir5wfj8clBoze2
lIAyZ1/l10L2wwp2KRpkPOUnuG8WKowVX2YSQDu4Eg8cyki7/MkV386UaegCqS982OqRSliZqELa
rFrcfSJi/KNsRWRk5dFJcVqL9+YTpiMRzadZflvvyrfTaGIL0GA4KrygYlfigq/coPes5SB3AvLe
GazbMp9Ot/hc2LkUvrBQT3iPbN0IWNXGrvS9ANHP2svDaRtiUPGDc264prpXdrSpVR8y47eMR5dw
OoOv61hIo3KVviPKAoU0JhyQBpC0xdzJEtz7vWeWv13562wVbqDswSddroGBO5p6kJl7eyZ96VkR
BLRONHITpbgZbT7sd+UdvBo5RM0wo9npZEhPTkAYGuDW7Mxl6LIEDQhkMYx5+9fxA1tWick7VCTK
F+v1FDXrO+TqkJFVUMrJqmIbaSLI52UWcQyTdce88OM/EQLH1I467zGnUZ6Nn7hO2NYJfI9YeK4t
f4y/z9cMbI4HtbfYEGfG6CdLo1CSVJxUsiQsVIQz01MvvX8cqV3v9752R+2spjKYI0llsKVKFFjQ
yvHhmKiUqvKVSjF7giUNTO+NdL6bdzOkH22iW0+K2tJ3a8IPvg+iNk0aW+MKOnwAkpB0lvPN8QPp
mAts43gEWifyTzeJ+KP1xid0c7AwZTxzryD3mjKow7a1Dpaj/ZCkfpyE9UKWKq7gNUq5RnTEZDg3
ESr2BBeDFthKwu+lT3C55qxYUHJEkps3rvlIifQbjMNIvOC2fWJo8GPSRrpx0lNQCLSCKJgWB689
89a8piKM4raEFlo5UvaXqQoXkqk2PJQvUFv2TdukIr4eDM75aPrehxUMno+72sROnUT84oZar6dy
YUC25iRGnmpaR3w4I/0ucnPKb/Fip6bNM/HWBXmf7CyrcvrhlL6XI8xOLgepnwOvSi4OGvrtIy7V
2ahCoPY1kn6zJdm8x9APG5c74gQL41ATkPFIFo0y17/icxaAx3oI0BYl/yEhe8HE69lDMEb6tTCc
M9eY+IoW4g2pK2sRl1ShfHVBgsg5XWtw1Oqo/IoWucQvMGDnxj4ljVG4gVSJOQVzT5Yy93LqboJL
aMF/yKGAkkLhdHG2KogCHCRcRSgqpYL1F6b6hm0U+lJhJmyOfmcnT8ogO8af98uu4pvYRGylK5xJ
UAEmkNuGDsjPx1R+Fq0EkDf8kDd1vpvFW9wAb8SOd/JJTmxA52QFyu/YOIv7ik8z5pYXme8ebims
GsLpGMNYLASdRUOGjfEYC7vUe+aFX93V+7MnSuGWEf1cRmpqq2ve8LADul4OajvgWbFWugfLouPD
u8iaocZONdLZOC+lTIpKCUxb33V+gmV9k59XsjccbgCVhMEQiKutn+lWw3whKdsHd93gVe2TkM4f
4zgvaHDjs15khpx5RJJmx9zT7pd2maKjc70QkiUxbgg6THm0+fmLAePSj6jRUvOW/IRVH6k55k9j
DDuYBm84bkPmuU1vff429wxVFkjY9Pd/3HxSmo9vkVbD8bt2ci5ntrriDlIKuyXTqk1WKUmnkKZv
owDhMy+53Jg+G2tLvxhKf0JZWH56BXHtenQ75RdEwBo2D+E+fzPC7SdKgLkV65hc2qqmFZJphb3H
SjM+M8qjO7d8IcCPXCEppiF3KRSFEiXB1ZoMashKMiCuo8x6M34zD72uJQzkBOmTGGsO/AZ5vfh3
HfpIDzh2BqsLaxdV/iA3WjGTfoW/TSujQOUac6rZhS+ERy+qIycqzDqifYIIqyCYQ0ENYajp38o1
XM24jSCk068taBk5Fhb8eTmF+QDyFB4OkNJtz7qc/AaMPLDodgMRIRO22giUbUgeT5sKzakQkhEA
IapO6RL+o4edD6Up4qYgdJJ3mMaleA2uye9or/W2xF2nZeqn/IXc6+g6jaOMZ5LacE6DFhlnhjFL
Zp4MgH4gi7CqwMxtZ39gzfDIFY0+D8lsbGHR9K8d5UTi3zeoL1s7zIqpgRjPWmwiJ5uGtxD3NJF6
yBfn7qXbdyyu2/vDdnEK5x9MgihLBS9bd3YlNemovMaxcQN2hlEqpvCs5axmj4m8d1KBIcRXgzt1
khhcBEAAJzWSplBbINp99Uaq4OJjfoonDqTU2IjuOTCRwFw/ymPM75OmXELRWqYkayui6cjr9aSz
BqJTevbMxwjrqMqg5DUtyvCtbnoke1b6Q1nonkEt3mC6mU5w9YAjnwSfvDiJXZ1nBon8HYJemreY
tNhSJIevV0H2x08VkIHmWq38E2/EyykTqaACTvzxO2RxJP5uaXJbuzA4NMcaU/PcGg+9ROcTI2td
sbpqp/c92izSNtNY0xuDmXeG+s2Ka90QQVw1yRJ9mlKNw+5+weg3ZPRRtwgMWc6p6F3WEcbdfLdY
hkm+fMzVyZiWL3mExFcvTOFIphEHnViKCk3b2h2y6EMXuPKej47uoy9bbze1VxgTbClWxB5xUlEz
7blrCskgM27aVXZyiR8be6D56c5EIrAOdah1EQvWzGDUcqTWYSJZWTsVHDhDvjXjdH9G9S26o6Ez
1Vbom50LvXpHHVCfIAp+E353xMO77QT9RrK/V+8qbLeN3E9iOSdyvy9EXLN/NyQsVKIvTUHJgUgE
uTtsLHa1oKnKncI6l1OyHhf9J5dPqIjvrItnlg3H/Dn+abZRbEaiSPdNBFmDRgWHu7CMuUq0QLV2
EIvR7saxpNiaCDEl30s66tDhKhajoXZCwEmCcHRnILTGTQmuEvUzrvemwq7a58Jo5sdcTktAAz4g
srIH8R2PwMohq+njno25YAY+7YSyNgCXOAIG7rVnCP+71BdW7wlI54ynUjdDYEblnwyG88BQzgOl
40KFQlxVLZ/8bXyQWeFcjkEaJJ0nACuY7aEMg/NKNjMiSHssLWChESyfA6Lvk2K7dewMFAxpgCh5
m0XSnk10m2l8dMYtbTy/A2EPRahzsgB4zghWQJ24Hrm7EUw49gZmu2Z8A/1BjNTJJRISDnP8weyp
YFVQwoB5n9EyP/M3cQlUFeDR2j8CbQrlOr99H/NVfrB4rPdc1585DPFg1AZv3iVW81XqOt6uCbQF
Wh8ardSUqZeDJoGIdaTiHAoLpPBJ+hjmYc1Jc1jWjlJnKps7OBxDW8edJXbkUHPKOpoz4C4snL7h
IWVtWLc4oY9gbZpnGrvYew6duYteC6aCNDgmwsVUC//htFekNCFS54egBvkStizi7TbjNqOtaazO
CUdH/Tbb9yqwe6MK4e1YqgbU5JbiqIwidxHJ3IZgDpbqcmggF+hmKpIOCAKc/Y4El6/uHU/mxdZv
bS2Oo5S82Oy9nu3XotD5+ViiXPIwBzxMlY3FWl5jltHVvtZaVeUlMQIA02RnBYU+53yly9nKFOKb
OZU6X5pn51pjIfcUxQPnSs4pa6CkZcGbIw9zuqE1YlvH9uu+Z+eN2jVHPfc82y+AEgqvjLXqK+YY
9YLDcaGFRTGUpI44hljiq1S9RiIy9U9JCNPymp3SLUcTg6RbsWVNFQWH7MUtph0m1QWX4oS96isr
OvbaLRCFI1Yz1PUXGZwbNfNPpzJM0tkvyALbxp/+/9OL7bhSsIKnHklL2x6OjE47tyinU2buPmno
i/kC0iCDOna7F8PaPt3i3sHWt1nQHp4Zr25AMTlld4ecQDPzMJecfW3AFyOrPRxr1SQTxnGHr1ST
htvdxDeygO7NQQCNGVB6SUhwEv9MUXxZFNNr87aAThUsXlpLpaVTrMgCNWRc9ARVRjm/FO6iEWbO
vd/DKygszZyB2lGuMbUvdvdJCivPSDANXXItFkLuU0mUtoS6GxUCDs8vHHKQG2Y94+Ydgvab6GXI
5u+CAMyOU0fLMmpMqRXKXf3Y2Dpncvp0yIacG/hmAs8Wym5sX/upsnfOD/6CbK4kcQL8BcmC6zhl
T7BY+0pMYRQnnu039v5WxHSFaL5k7lbY8O3pnW8XqVU76xg2nyki5CqhGTdqSC2HWbSYFHkUnf7N
KiZAl2dYUhaxhGUZSRxObLMJI1v4Qn1B5TwLI72gRGhZkienUscRKy4I5zpFAV046pFaxVrfXjBa
E6JlT4s8W1wJ0s9UJ7+aQV+E1IKFf5WXAwsmuA4U7hRjt2UYj1hoPZFPCWCp96HKEhw5leTC4TKW
8MMbraVlvTHMLHpYmZ+fXMSX0B3+jQ50iJPdGVzpzK8RQU47EU7P2og/CFoSRTvQ2xp/OTFIo3fu
rAL6I/yQSu0T+M69+aLOJpBx4nfdcCil7aZxAP6tCBlEYsUdcbCUD7lH+5Pov2DB/zgQgI6qARji
mmWCSpLXK/r/+LfNaGcOX3PcPy3UCSMRgx47VWnHoehrY+mSzc+947/rqFx+29aMyVStaSUi3dK/
AQdNOG+HaGpkhLb50VinJCHzzb+wdmjo1w21zVMAusnTcGM04i8fFSfJ70yK4IxDFSQ2xjjJw2nI
mhYJBwFbT5NG79G5dRGr8N2xVZqkh51PtXVidRIU0xx+g2r3eGfVfw0n7EDRvJaVeI11xQr5M0L1
GLAnQ481BRkMlGRlR8TveOpLrBQmfyJY6IjTPkHSv2VCVgmD0kAYRRSHKjrtqBz5IeleqRXgtLKy
YkMofQRsr1im+EtgpJTR4tpgE9QgdnIt/yTerypcK/K8JTQatPMAAX6HJkBQ+DOktvqsK5l5/YpV
6rWcS/1kh0XWyH4bmZjsxsuLy35jDmLsExVyLs3nSPp2xU3mJZaCI4D8ZzAYKIy+Mzblf+T9TcRg
nIANRrd0zgETItHh0ih07HjO1WDLrW2EpIC22RhZ8cEuaQSWasVTbQfvN3YgaoshWFSt5bWTJc6k
Pc1UYciK3/rgNP1lqs90vhRZXoa8Ks3voqocPhcAdBTbqwAkCKWIyNCJUNJM1GGhb8JPqH9Ni6S5
b8DRWQ0PNl2dOSfBxsBPzVgEqZLTUGj3jnacPaKt3sjGqQtCHAZirViOXZNEZ7QX4klk/ckCB5bm
icQC5nydWQAIBr2yIXA1lBs5si1lsFJIReG8SuG81IcJhiXnptXmCHzF+kfVgR8ZJtY3knYhnmkP
2A+l6WaBeil00leQL/E6ZMjXFIkan4HsCIIX8Kond1HVCZxI8r0dY8/UQu/5o9UkRrS1X1btBV3o
b8aQ2oT3x610Y51tIMneNWcRBw8yZ+C9CflGA/DuBgGf64ISr14hfQjcLzdpbntvUiOm4kIRwFMZ
/bUashZ8o7cYojdZqsSjJrA66NvFTfOexW6gyE0/78knKOyBhrO5Ycr0Gq4UP0Ezmke+o1XGDbEL
yODPDjYHMjcccAzXgoo1ohbsG5qS3kH/XTAB1+1JGxIVaZN443TRjQkV4RmgWfM/FkvX594+25Ea
mUPrJnOZd230ir2jU0N1iueRVcWAbM4hQ0uDgAbofz5ousZ/yKig0lny6A2QDT8RjHOH1CemSSz4
TKTSiOvjT89be7s/ji1A7i1MnBqLxN+FjaVAdXap3bCMtYms90ZoKOGItxQ05kCuDVrnW5KeoiEK
kVqC/V+Bznnh6/biOB/U4tpWsjyS8xQMJbxsg6m/CFP55BJtF4Dv4zqHK8DLzuUYJSgJW1hbcUDS
NCvBTutQ0V7pTxlB1g8dWH3e9I28H7+1a+ktpG7o+Z/shdxM/+W1vrnIkqgRO6RZQu9cnPom9a9l
LBU2WffkUCaNMC1MG6sOxQh213JR9T/IsOYNtcRNMAfvlBtXezeVKZFsSZGys6n2B1EnT8EaROqg
CrTY6kFNEQFa46vx43fDc936ZI69yTxTQTBxsfC9O8UY1MJDTvmP68HzUsTHrY6Pz1L8bggAJ7OX
9g9iAlaz5D4wPlsevrGog2j7/26uuY1BN96i16LHc9HR9ui9fOCDSFdVl6gJ5k/Wt5uwELF/ioL2
Kb34EbSmTQnatJgT0h2f9JG8sJbmpAGN4jLYhg255orTWh+HvhydDGN7WigUWjp51f5p42H0TgI8
+Ij/w9Y+7xl4KMWSocTIT2+XaAWb+0OOHPuFiwuWu/t7BsGpudkWaKIpvv6FhOb+kzLbCiTo1Xz2
X801V0HoUoisrohd1ogxVTFrgmmDl9qK2y6R7au8d7mDWX+d+4lc74rMpcoRYfkcjh15gAZD82Br
aB7gzvwQ/PJgYKIjLePdJgYq8M6ODlUlLodNVawsQix/3Crg45PQCaSG4B0cob96i8rhkAVUMrvu
dc9oeG68NQnnHr/yW17WLHZGiALrtUYlE4eMFb4E255rT/RKlBGLbT2HfCEXP/RlvWGGJ7FyyGEu
eK9vjXFQenn5MtNmgBzI+oNWpbKqnSC/SB/YppX6BIgTPdG9YYXLEQ7MBmSwLrLI7O2tdAzKhPTK
Vu2b/94xOvK4eJuXmh2iTKmyNbT2ikOFnaXjmTrKk/IzwTCnbVaOLE+Vw/40Msvxanjrt2vXFNKF
39+JcetQW6nAV6xU7XLLOdsKyTTmgk+FOS2RuDR2yOkYuhbTTHpHBXJRdEJqvbkw3ZqRLwdNb93F
dWU+l8zkIbApdslCoIM8dQlgNrD3hS0m5P7wX3piH7XsbABqPhDHVyJUJ5V7yOH1X4Byp8fVKIBD
/EIEr+Ej6Jop9BIDjOj5pYqWL5ueOGwYfjvxTiR4XY08vpu1JvnfiRMPAtqOpB9yxWA6zcMNjAdv
t03BbcQPdUod2LK6aCdDwnHTTgXgxRHovLJkn6EKqWM3AcK3XVrOCV3u8HB9w2FIGPzBg/M83Jlt
lAKC4QYfgeDTb+eXthzWuYqO2URbPXGLEaEsfEQduA58U9sqZZt6PGv9SfL8+MIX2RC1pd3d4UYs
uDb/LEqoiQzg50gjBG022XL1n3FwyMVJFpieyejnXb41ALOvnCvITGiMdiL/6EvmN+fSiLwlAoSM
KsNZMDZA5lE6vEMfcKeU2Towlp4ta6azuFX179Epk5EzTuNolANKyLu3Y9YyV8hM/y82iJPuPtkw
NuwZI6EUpV1WDxa9Bq1fCtesmnATVkpgR3O0aMjOGrNymYpfL456CM0Jexm1lsEoHS54DEVpPZvt
e2Z5YVonZJ1gkHsnz5ZdSG0zylsa5Uf2gZaQJGIkKpdp3v+f2PKeuwYPXLaKJr/5QZHNP7b7vSw4
S5S1F10tPCjoHF7muWIv1MeomiIMUhdqGWHhiXngVGkjZFSjZzDwy4rRDBK3LEOEvgGMVdYqXCbH
CednxrB/1E+vpWxMzpRRMEdCBpAncV/CerFnCvQvpYvGuiLdZY0ZdvYEkwVnATz5aHqs61NTv607
qX0ONfkYB3jlvT4scGrJxSymmnSUkeW6mXuO6WgdAtvihkapym7A2PLj9jX7wFbMecFbOsEssaO4
9o2qAaPrLm3+V7CavQNmNP9f9NJEmCoDLczXApm5pC66FsgyAKZZfNDLtwdS4nqmUXKd6+SQ/AxP
SIlcGOxM1ZFCF58wBksEEOkpTpIHDXdsVxdEpql4dElWH53gogfPCCd/vZ4Nq8A6hE4LVhn5NuDd
8KmhS3q7aY6dAedvLQbSO1jYwPlwJG/d/1HBM+Nkz27zKUtDVqXukVbuoHseASE/AmbhuiD288bY
qtzPKtJx0WktRadewn+mNJS7DFNJyO+gTbgwtmy+uO0Wk4S7JWmf1q3wVwytH3DAKGu0SXk0leOy
OmjEaTzbbzRJcVqlyA142SHA1HMAkH76iMmN8hv9OTh52wAsLaTgvO/CL4umYtDe9ka19CM1lLPP
r1kHti+rKRFvzIaIrswCtQ1WxU12JsU+feAwxCbNvGLSPkz+IrDuOCrCcJKPURKoJkfcbUU+rV8y
Ed3bgHRfm4WuPPWFrAC0pBtP2SDpEW5SmUZ062yN/g7y6bxEsE3/zVyaoMYTLy/PrBAyyf2CrWg5
UFwfc2EXztk/m0twf3+4Zfw0X8eYoczhJSl9AB30Gvw2/gQBFfpQkPiEEtgtuGb4mVcZNvCeKDnw
dDnnE9PXGzLYQ0Kx2+wttZasuLJt6mbkn7zqSjlW3V5GOhgaaUJBPgtkTeyDB3NIMz3t/vpgNRFe
deLrDpxv5ooRnZ2gIxRqjsQ0GMXVdZaP4VQsP+BoDE1hID6DVOxc2RT90K0erVcy6BH43f9m7Kha
RtKHELTsFFZVySdmmQWlU4wTi9kSp/1zfYe2cWLpDHYipr4HRbmmvk0BwfFXyrCbOwTrwWZXAMbU
hYrphj8IKZKm9jz6PeN1o/JRRSd2e6D3ov6MkV/8J23RXXpgEeSZt5EwVQRlBrg1aJ/Q45rt4O1J
xgKJjwBN/u7XOs+WV3jGA6Hckcsx0ySiYlhppTsC8jgECKUNW5s9BJTHzV+W4GRAGyr1iSRnNIBx
TPFS1US7LtiAuWOMMvC1iHwrie2bAmqfkZYINHIauobHHP3eTuaHHCcjZ7alwVDWNJvtbaXZ/TDa
G4pQnO1h0N/up+jM1Otvrm4tShS92LbvAz4UWz0Uzg0F/EWwaxvXEvn2tYW79xqbQ+zgkmg3LZ52
ZLkjseCqUV7JyyqSSnrA42bPdsj4nlRd8/1mxMYfq+NyPtQkyrOb1hwc4w1QmZlJS8RECT9ubSpZ
JBGqKauKgf4pXFdbcycQVJIe15U4Ixl9XgG2IJFHcdkf47adtGPSa4IGBPNOxx9LDgaBIAAvyy/R
VOj8+ZCZFFkeqHFPhTqgkk6uwWeDXB5wpSrLCS4p5CWw50oOcq1J+a7oZ5brjzTMSD1209wXXUui
gXLJrklvkWwb/gdMXS5qQCIoZhTTbevwktRc1LLsmBR7TB98dYr6CeplRWbn7AEaPPak4hG84l3U
/JwcKxD05JG50T9YTFB1tKmETVWBJj3c8eE9jLz0kfudG3yiULgTxzNMwp/nnoUuIbXwpXUNPgCE
FzFsH+5SSzwb06RUORRqd5R03sLq+crdaLZ98HM+E+1QdiYh5U60EsROp4L5CO8iAu9DsR5NO627
6mq/vq0xNEdPZqJHBWHzW/pE+Zmr00906lfCNnhO3G8dyp4nfHE9pEXu3Rq9rMm0nLgUmwILlgSp
Oltj2bRZr0OsmbwigWV6ft2WW5EUCQZXtvnInYQEXKXGR2EdlCzcgu2yByVSTiItufTC115wsdVO
9mjTdk/DmOCYnVhFH8U4Gn9pVhvyHV3eg7Z3gPSS0lsISKJZrZJCz6uwCcxGUz6EQ8euXcrs2fW9
+M792bnObY4aziiY+fyR81eKdNmxJwrhvnc1FGpenttRv1zZvY3al7jUJVLtSrNIgRwLghGznCTM
oZzXDDsJSzImb44ps9uilQ+QFvk+cZTn6MbjJA+dZi87MJKZzwr2zquOCW7tx2R4+bWFS1W9XwXc
DrGJ9pgxMJmTiuzFWCSlu/wOmcnDR2Zo45hTPzVfpR8sDY6bkxhMTvix1pdtF7WVH7nlrYS0c1CI
n9mFkiOjjGJpsZv/dUlYTHSgO1U+BoymrrsBrwDa883Sr8WQTjPEfyBXlZ83SGzYXIexwomhYSPK
8pEBlO3frFrXsHN+xibOSlRuVUDZhye6TdFFckTCWbEzqrxJT1SrPtiZSSB+u7sjINu7+bl+hIoD
yRSVI4BPo7KTgGWwkNHPtBsuZAy8ZvdKqnlvTwJUZCFMtE1i0ylWTlZz5Vo/et4bMXT2jrd7APuV
jtaQ80/YPk73C1FCGQVd51mq9VETY4rVOmQlKcpfmWAQK5Tr1XqnZOLnoWiajf1qguq/GIOci2pt
TTsN/K+VphztCrbaRHoV+SXzWc/Cebpf76RQXDsz4dOWRECkUdKbQaDj0HLfonXiH/MzgW2H7EOw
W/c/RlFQCnQ6pLEdrN05lKmLPpjzqx7valqzZ3bR4s03uyIjJpp/GPHLm9bWJdp1lG6Pd/DozSjx
o7vQyGDg6tcF1Big/gLqSVzPhUf/xKE3tf5MrTLd1TAdN+RHlr9MpfoEgSl1cC0JhJSLCjEWLBSR
Axz8pTL7Sc2GhvAbnEX43maHq/uOkZZER9Je1g51qI8a5Q7O+G/fRUqR2JOJozpOOIvShPRire7r
y79bDY+vSYyUVVIGhqGzpER/n3FHJ7GLQB4WJ4GrbAgq6B6dUPlCH6QWUyTb3vIqV2tmQYJLRax2
RoYCZX4i62yvJeChga9qtjGjQCRpqdVVB516P4w1aM2m+tCuXip4yKieSff0XBVyaNeDt2BCp8JI
JVwFQ59w4XM3i/O5knN3xX4vMIi81NCZYr5IsL7Te0oJ0Tz+e2s+00b88PwnPrGHnO57P8Eicfdy
lQ13g9ENquuTlAm+ZbIRdZgE0YYfvFtI5kIUlPTb9sC60TSLQhfXE5KfidUVNLZjj0KWBL6Rv5Sh
2LvEEZsFZIO56dcoFux8E/bfxl6G+HV6v2SkWf1zJnNhAzsHBOz7GsIKVWocO13oNfGABhy2JB0P
EE804WqhPzknbANDdLSUY41KlqIZGyDfUzfPMsDUIz/jQRoXCtMKZhX9mlOnDh29Gz+6saKf+omL
t3ElIQt4pkBHaWi9pV+g9mkqObJFB4n0TYC8lyLokk3OedE30dyfEwKRsiisjfKhppVUwLVPoIJk
U4caYpvhqQ3/BJQZuVAjnJC08KZ3jrEvHvW1KB3VJMrNDSOgV9reiSdsRBWc0oUNI29i/UmLHXIT
SrLiOHRXCFWtr5+0UfzP2UFl3gUoaA7DxQcciz/LjdBbMYTtRie7LFlImYF/WiDZ2lBiZ5/lKpLn
Cnwe0ywOiOJXJEAdlZz0TC+babYnvVI50lDqckXAJmqfJ8aWavINjHBc1ygPdDvSSZ3tx8K8oJ8q
tRFIC8Bmgori5nVI5On7+eNpzAS5UBZML5a3T9UutLQNqVIr/cCM2zJMnDIpqXSEkvCNGEROFoj0
PVOPtnSAltkejfE6AD9XeZLnktcGGCg1HHey/K1/qlwomfFKbnN1A4mD/y4ULkqCndb4DCrLKXpI
top0wlJ8BLbmN0MqMKU64aLs/VDLIq+vo/fGCyqsAJn8eqJLYZthxW1U8x4Ky+aH32Ihm5ufmskj
2HJYaJe/7N/u6AqcFrkBYgi4tzbxRIrCQX4SQdMEZbBhBws3Vf0k3iLHy1KN+zbHI7pOF7GVs4lk
fYA1b3321SQOfLM7gHj7zTsFWp4dq3OClgP5EJn2BnrpfvBPH7RpS5dB2U+VVnXg7YgEgFCXss7S
xw79mVp5bzCOYRImc+9aXmj1Wgy6X5i7E3WJPI/Mhsaw7ClQYaGgqrtD4oyA5yurscsofHSgmyrP
aUzTnTMqwnq7hWeQeItZW769f6c0Za+E8mycRska/a1sNPRRYVellHQF9VwO5zLRO2yWPrerZsmr
XEGwqZIlj0onZyuAqpsyZ4nbzHCfC1jx11O5SsT7O4s5zXqNwpxkuBBxKRr+XfywpbcPlyLROYYJ
W+xKO3Sgif3R4XT3GaUj7DcPtIOp5tDbNRbUq4kseWQyP0pX8w6ZQszbc8axMaEKSY5rDkoPpGZJ
l/xFFP5TL43v+pd+qHMnELbaYBVonCeaAR4TfohiUXN3l1HCf11A/QEu7snV1pdcF9GXe+6MMu+A
OUxYb77f59WWnLoeVVyu1GYDnHby5NifEFVgoA7+hv16V4qhUdrAXbZlPZvaALa0dbNcebukGa5L
xEv2QdJAi+50MXxRZmWeErk7Ekya8+Uqu+6TGmU651FWMcttfg1qLGiliKF9YzDIPSLLt7ppybjE
edhgPEb6zZaxErGO3DBrfaBu/q/K67SIzIhe9MJoVB3ud00p8m3HjvyU2OA61W37PrVTZXCtxBBS
UIm8rKRHCQq8Q7iYHpCoc+MNGspO+BpCXX7PpqWrrPIx1wNbWOY0rrjYxXUJS/Yk29/TUe8hWO7U
Yqg9wQoBcDHDNoojqvsI+Bj8spBNN4RgKs4h/YHeFm6iXr5HuryFg9h+q6GyJURi93w+snIiLZIM
GeDtTs6VxZQ3fvX4jBtwRXVvsiSQ6G2yZeqAJRoXYvxq7QduVvHQ+0mgrTE4yvcY0ZPRtGLjor2t
VzO6HfbrhYzIEFJ3dJwICZPGeyGPqKV8RYPYTbFrP+yUh9YhGzo4thF4FIXrDT7RaIdQ47i1w5f1
3kFMT8r2nhQ+yPjyig7YjcpGT+dBkt9+7xqyoliZOA253DVQ1soEE5HlprUyH8C+EzD+uIC488oW
p/KGULyzbWTZcgCMFWgoKqOwS/Y/hA8ELhOkf/gP3wlW51ITtggFj0cJuQ427ojVkqQbK0JWPzPu
Owgjc3CYwUs/FgW9yZaX2tMEKXBEzNFYszN9jTIsE0SkgM8bVUK1fJCUSPJpZ5lLSa6YIVhXkpGu
4Fj/YgkwYDyTRQOcExCqLFomym/k5gGxQnvPTTQFYywHbkoSGvsVgLyBq9xEe2SpoPLe0/nq/yJB
1ei/kzzfeok8A+s0wMBXiiu7SJMF5RNuuzHwKrfuvOGYmPm9GfpaxM+ZZiKjEfidVBW+ijskkpoo
nIe7woFH7YBS1x6YIxawsmG4lqSKlc/5oC2qNmWU6tSI24QflVKXJ6sieUhcucmWUqQqO51oX0wy
qsl+YHubcC6gLE0PfFduy8OCItUZ+IrtXLTbcc/LPiDdVF7RmYDdDLf2X42ONotW+4VuV1s/lFbm
jAAvi78PpRYbd2XDsss402PSfVj+dNBO3+UzXKw1vyZOjtTo82dQ9dCcrhWYzH9Y/ko7vEu06fQq
leOVgRDVqDAulCRUCAJQEp7/zN4bSqTFi0EOjlUq9WOOgWEEX1lZejg08I//mS1MaVhaZHinPJN2
UIKzqQeRR/j0to6BUl30EqRji/ZiXwMnbOUKEAWbnzpyVRY7MrJWNHklLxnoZ9hnUpMAg3ypBJX4
5yy4t8KtLhg3JebSGTj1aOJQCyjL9Bg0rbplrWJJGhZ9EijrtEt3+7oCbPMEpSp8w1AAdx1KVPVt
TIAfpcmuX+6XqDXd/P0iGg5XIMygzWzDBsR+jLGOzhHmASgmnt//kz4qzNa4KsoTVKX7+lrtz+QQ
l0HQU1RThRNp1eEHQSXnLZayD69wWz+px25CdUbfNhZm1hW1yCDopinfc00tU5Pok2SPK/KXNwMC
60Sh/H6ZN5Sn9viZ+8eA90k2NSMfocbDOjD35YGHq3EHF9KFuoAkZJfVK8MExakiwvq52ziKLg+P
opvSkX11S6EvNq+vOrcBXBRzfVwUu1WmGW5FofsICXMhk+D4MYP6lpYwCtT9elmDS1BmOJpeOjb8
WvYSi6473GvdYcBRatTnhkzvG/SIUHEIS1HZ3W4uZadsaSMIr0G8DCak3r/bFP+sTGPDpEObggfS
deZcsDzdvIBp8Lx2qGVhyDS00H2zoPtCpc5YlexiaCe+8dyovQfUK3VlG/8ysbc2TwudyWxE2T38
te2p3RIpjkc+WyOm/9Z3hY1BbLrKrg+ZV1NOryBraJeGMmjIEzH55xDXTkDPMKyR1BUiVL1VBaqG
E197AMC/7nB25iC1zaaJlf718mcn9hKi0nOPegrCCa3BdtkIjHWwU4VXpB2owoxCVNhS1hZd31Yb
Nn0DX0EWZBZ5wHphbLgknmXvbZSUO+/9xbohJZOQ1aoqGVkixq+eu2Wvgv6qLG4zhmoVfWAtzXcb
k/y8eL82dX5rWCJv7L1spwkBxbV4XLuHh/7M0Bt6rfTfMa7610PFVQja50QQds4LL9TNfmseozEA
g46cRYK3V4QpBw3ja1/yu4SAaWD1NwpKplq1m+8vG9srKdY2zOCRUKRAMOF1vgiVUQFyjas9idL9
9QUlAGPea2UcDr3EsKTqYU5i4TRp6oRwJcWtcbbFo6pVOE7YRbfw6suXeY2oJRT8jeeymE+B+4KI
K8QwYiNf9KpYi9nQYfvzcl+aMpUtwpX7MCkipd5H0tRy/W33Y4D4vMh6vwz9KwR+lGm8BS+6xuzV
fNnSegw6TOjVKSMzB+zLTUCVmEcPwdOb12lX5mc/KlDQhhWiSY9+4Dt++bReTzM9P1tDey46eBjz
xmTGw3u2ilKizaj07dcQuilUypBjin65C6nRd0jq3S9S5RL1apkyOxoLAh6OebjSy/pr6XKStaZd
y8BylA/ggXvAfl0Y09PAvCvOF/MeEnTJeow7aoJo+vP70PenYlApn9b9G7YZqIfssRb58J8SH6PA
2iz5EF8YtDLUUoL9KZjhVyvqK9WCIDgGXIhppzy3Rj0+Ug4DbbvxVhO0RHwG96LAKWPDgowPZDvK
RoOv7/8bVXXzIq6swESoqD5uyPYXguo5kaoVl/ynvxmaARMtoL2xh2x32QGLq7r2ufLEkWX6ugtc
gGcKYJIXwAMpmC8DTqed543V2vuWbCvV64DBI+S5iIBmcvE/s4yA8kFkfToZQ3foOK1LxsrtpMiA
fIrZhp4BUykqg/eGvk5zZqiuYGwN+0Zm/DnHvAvedGCgWy8EDBh5Tri3YO8ZM8I9Q3sWsXytOdhf
Wv0JOCRtKi9WldjhGl1vdheH5wH9frClomC8iJe7JnawYSGBXOGRYl311rKHDNrxMcHTCCglOdk8
exX2zNShIz+wJmUzjT3VOHjhtTmQpVEOMFSoG7Hdj0YKRA8+Kf1gC6d2lRmAVzlY5eKf/OVd5JEI
2/lwwK23p3A5dmMno0nXwnxkm2yv0Fk/SSCXLjymcMdTtoRU+xMWvP9aYSW5dKXDMR5dlJIhHHeD
PgbDuwhIfbkcn6Aw47DSDx1GCTgEwRNqKxBEQgJjLbgdT53CCZmLnuktFMB80yCPt8V0JSv+GufI
LCCJqCc6SjztbM0K4SP2yioLT0nENIpL6QuCTKhDlgGg01IImRdaqEmZVMI2dFXifdoLsnmgUzNR
WVOys6e3PUzoh7VVBo1NADr3iZNg9Kxa9IRK9dPQ0yASnPIwnov9H8ADOpXFK5Hw8JRyQvJURfYB
Aw4RTICD8M8g9/Rv3M/IzPIFsRMRYnPeV8Q9JlOJBsgefLhNJg7b9mOka/gGCpgwrhfeAhVxDn0a
KUEGDnh/PXq3xhAJXaU4M/qyU9jOqyeoDVuWQJf0HWCrFbOGDE3cYjZhdW2b86Um0zLoowsaT9vH
B2Iq6CRfpqowVf//vYpm/dT+kgAd84dbLfeB3QYBtsPrbkKmPnpBSzmWuR/BcbM5rzRCnK2AXi47
aLU4IKuKdAjUo5XZRXNB9qfS+6WyF97EznBO+88vgG8EPW4WOpWZnCz8GxeXh0Zdhl2m+PsivjqB
Rs6RuaxjUwGMAsjbl/CiHUFI3cSqNUcir9cgYfd92mlW+c0ELBTWjM2JYud3qfqhgdzyoSA9S2qQ
tC9wvnC12k0FGNIRhW4iUQfM1UJTD1fFYlG6o4yWNUcfOf4ZZWwyjDoso40Pp3C+K0tb+27uotgQ
Rmc4MQe3vVTGh0SxQDLX5ua0imA9486eS9EzkwyBvUnp2Jz96V+je+KzJ2pUvs5F8/pXrYh1sndz
zrS/4pZY75tu6TAx7XXmM/WCm0z9gJhwH2UZFuM78Hcx85kCjh1eT8XUhcvJbp9Ccgva+HWrbZ/0
yKw9DdaNIU0qVNnggK9pj+wc/I6P7fIMtfBB9PaUH+R7+Ju/tLzMVE0oOgVyeS0kfAkBclYUAza7
UvXOpWSojf7PS+IE5upugCTlYkEVq4A+K/Fqaqq8eDp4acP7Q5aXBWg52X6G9F4a0SN0edtm/Du0
f9rHRyqC9Whrg4RAUNzE2edJUs2DvPjs2ShGRjURjK6wl61Tr28KrEzhgnWhzzJGt+xVMjS/60OB
EHwh5w+mzPvpVrhU/zzdeG/QBRh55hhbOiHjZMyem0Dfy71RVQODHIBEFbxLUHqXxd6NE4YemvzV
u58txYbwk6GQ2cFi82X9PQfs3ivdrhokEL7VD2GGDJkDLXlqmuVY76JJwpoJUz6rsYYkS3wpbEgQ
3zMQalVUPJwKkOU5jUI2x9oR3IfhdT0Ooy0Vw3PjwWfaosSzmec+S3I521Hv2IP8lDJdkab/GZcE
Wle8sCc9p4nF9b349qJw4tGgFDbbxszfEYrZEw+B2zK2/zFErhWDBRGrLvVvcwP4ECrpc6xUY76Q
tJzxThVVYIV8htzYoN6OA+eiZBWSP1r3SOllCtAyIrufOgBO8weMJ+QOLUhW/3f12SpaxFStu7h0
08sCyW757lGZZHaL/KEVRmZ8XW3Kv6rwcqW5EeOclw+j7/CRjF7YyESgPhiVPcIs1tuV12big91w
qSFluXHodlJKDy9cSXCe64nhaHkwuIrPSFRjqIUUrZkyRk0jkZy+YtWerr88b1ndH7vuQISHqgIJ
M9am4g0UsGYdWuO6ole2Iog9VcAz3P0AkZgjommwjFX1Ny1zzg1z9s7bPJCciJeyccRW18M0X4t9
kw0VvFz0DUvvB0hBDQYgHBmfaGZFrBYj7RimBV/QHYDia6asdfaiqJNDt2Y9Llz/bBxZIxmtS9HN
xBEy2EetQTcDv910GhpVMqI0Y6eXAQAwwKTtnBUrA69p99ts3+kTdj8nrQohvYeQSEQ7QHVONT+2
CPoMphDA5zQuj+yoSBd8+azpjWf+2lUcBCxV8P/9OKVj0U1W9dMB7uwkd9mUFU3J00m117DFuFt6
n1HllhTSvEfyV6syUy7x2/kHyZ/d5MDO2pPWQuHmeq0dkqasjpsxvkVHl7/pG/NFFwBi3X8JTSkT
y2yIpFkzfh2n1W+BeBEcus4Qzqel+kARa8ce44xBn+S7/d8zVpDFh5VYej0wvZh/M5+lBVlNXtAE
b+MFxxGQgOgsktZ6aZxh59tzCJPunKmdDFI1m4p/d9u9sM1ckq+Jpgjzry3W+Kt4TqJPXGHuGX98
GS9BCmL+lQEBDUqqYtfPgQ78Re7ceDpzkRfZTOR+Yt+BSW9Ug3ffqJ0wPtegOTRd0qkX7G71J+1C
VebrFLvPuy2vpN6JAWPhOIfIEOUCV88rGH6S1gJCi07rth7M2eXBSHrXU2smrIhcoGx/Qh5HlGL4
AqHxiHWTqtG+Xbht4pc2G7pnbrnKj73DDeGAw6/J80z4YwR7B2sHLL5JHvBoFwGSs9UoIoLGazLc
fTV2ou97RkAOKei4NmiKyX0+hau0GvIluaNl0X/IdyAGSWa5C2F84a3u6CO8UgP8XU3HKTbhm/Zu
4VQVXXTB+9iIzlHJl5R9WiJ7H6I+1feH6onZv1fO6UyDjJlvpwelZTJDaP8EGtKFzdIttTJwtfXh
/mhh7OtHZWW3ivfYOllgiFZYKOPrmWqGTJedIF5tLF3EMgSff+dPnu4qKZBTEwb/Xp9qtFOsDdW9
IYKv08b+/8fxWfMgyhSHFTwd2JGYs8jT2Zprd+xA3TBM+hf5ZDRHjcxJ3A09bIXXageGVAWw77g2
2B4M/XeE3kLsSlP7N35YmzfcmyrFrdYGHZ83gGF6xDIXmAUDZq5f1fkk5HaeTa9YW8DyV4qk7mIp
X1AqfR4HQcmoJf6pUaPFpD6aOvzj1Z3vaacHH4/WoZ4nzxXh895fBr5O2H6mATujN6HszBhox04k
/YXSMZHkl6qJAWnkZ1NftGk7S2MphDiU0ls46RTCppnB+B6I0Jb+wM2FyCTT+uhZFHgm0tY57ziK
4T1KNsrKePnBsUE7sQ+0w6UEsye05pgfJ1kOHbxCwIqYTKISnhoBAZ4+XlP9pU51WGk4K6A3s5IZ
SEdy4eC3zB0YPNgUiN4zl2lBI6vKMXZYSTCwC2yrViTwnhF8wqeVVXa+cxEGs7JdEGuXug9jCayM
6p0IJCyezMjZ2HR4rPiG6mDrmaFhC93jeujry2P2cs213FdJYfSEacd1A8Sg6yiKkUjT/cJ1AaZs
CRQ5PFS9REJg5U2TPvLGpTKI93Ybwv0EpdDibDxRTPk5ZWVao2jXlX9brtzfAMCuduSOM7rppw/4
3FV5YM+hlf2llXk7dMstABCldcQ9JZazMMX2CTUgITe/vWxI1qkNbBeY2vpig2AqcsQwDwlMCDZ/
BMwBxDX3TnYxZEwBT5IacKjnYAQrphVhPYIIaSH5MryIOAoTxv3y63EqnmF+e4OH12hS/p1KuK1X
HdzZjtrBg6j7lmPbnTxy6Wf1gEZj1vi3Uy5mE7pl1s/aRiQwRkoQBBtVptJhuLFAmpon/xzNI/DP
YscGRTXpTYUvHK41TegnegSq/audQgtHWm4GICv0n7dvoXu5+GcBkAJN+ZNFGMgEmepUv6CoOFUm
Cl7KH7nclUDQuYyJv5c6Cse154z66ilgCHLdlGf1n2cLA1rIY3HBt1TFnF9OVIkVpaC5DMCzpWt7
5ga6NEIhVTUiFdt7EQQ1PmEeD03W9jhXnI+TgUMgyfb3JQJUPTktIPyl5gw0I4K+KctmRHq5MBle
JdBxH1fBAXzGq5Q3DFRNKQS5Vk4RIlWTmwbwJyNfZcw5oeFLVBeAXoxDvSVmm7+tlHyRVerf1rcN
EH1zYu1pkLoaBsC7y1xMwlaR62G28SfOEXg4kcyAjJIStSBpLg1mSNWv8Qc7nOK0MsnoRxLXllzS
QLfJ2ksf758d0a5woO33V221EVsKzy0rsnKjiP6rB34LqWmJbVX2f9lI/ZAAprU3pl55sJvaPpID
Ht1PkKf8sfxGHt1RZMp7YR75dbvCCTDjEb+YTmKaUrB4Cg10LCORz233O8BtJuP0tdMDJmBBzLBT
49vBIO/LOY/IzWriExw3lHnU633f3n8LXgz9yQBttiRP7b6nJGQZaQqCliQhccBkK03PZLrbTIYl
aRWS+XiHIOeDWOZogi1RoFNdGeNgJzo15Q0sB7yTVVG6CsMFcNJs07XmabIW1RD7JUodXpM18UeD
38hmArd1lDrkFc9AZAJkeV9c3O4XdlLBVd1dPmIKW8KXYBs0+CvsTzsT31zwgvY8CpAzau9nx4qC
QRxs56VXYRkYTQb1i/c7ooOWGYmaQRovCrhx3XUALHxOf/wfx3UcAGprWmc3Xx5qKsbOZyom09Gk
Sv4YknYfcxSSIvodTuw3RZ4glmbfb2FXYmakBGdi8+RT1mz4diyP3g2Z/vJ1hwO82hRgVCN5Gr34
y1BXYj/kmThTWokrMTPIKok4lfGWruvV157hPIgy2GvlfQr0vaw0xPukzOImwoBXMfdInryCe9c3
/jHBKNSirWWJHv9mDYdCOMsnIeLTW6lcYCyrL7rLBiB/Pb2v0V73ciJ6gSF3PaMmUVTFTLRbmaCZ
YkfxRvePjtfeZXFk4KDiFvCPfRc1iFIabWeYmF5J97sjAHacExyj9nnO2qFaVvdS36PVXqZhQ4X/
S4m1W4nUKTXmrZZw+j0t5LgvV+WU1AX2HdMKGWCvciOxBVCB32AwtT7qi3nwYX9wXt7/ThahcO+G
C+KC92swW0p/wQLQtWQRSQdncD9fsvGRXctGlaFwQkKpo98OlwUz/TgpII/+AZb/5BiAIYpREaDT
+EH4I3j9n0b5mzIoLIoEqXM3ZX1EQp+YxXGK/f2InhaR7rRy55awHYxGvvMp3D8lJ4Nsl2mvLVmo
VwG/6MOvN+toZqDWsnCa82Hm93N5Z0We0GDm1vhMcClDiHnDkue+VUwqShmvjrlV9DsbE01ExW1q
LpyX3RNqLcnbCKLIOekop+TkVotOUPVdU2LDVa946wFEaSgsesBhUy2FVIbDQNCCh0bOcKDm/HzP
AMvJM1NSkc1YL1NTztF8f1rYzekXz10vQtrep7qz42v/J2CZKY5bKVWFBAugYj8NpzUqUJee+Wa4
vSTAGIAQ8NbWv9e6pMMJIBZZtmEAT2CzvPn0azCRKseh7Q7DaM8PV0uhmw7zUYrSVxmVrndKvdsT
EmDS1XUtgz4uqGtHacw7uYGWxCKpZY3QvOvzcjHPiCVPkbXA8b8l2Ck/PWJFZ/KwehEEBJSAutV2
J9UZ6t90FlOQ6ChprkQ3UeFNZxSkYjm7cF542xeRUBWLddKncfecxw5N5nKBYNwEh9kolDK2nk6b
0osRFiREUWoZW0ejsm3pYN8LThaGAzkYcvypEtUPVBzNuJzqD9/Mof/B7uux8wSonIcyfklEwZ/n
lSrvs1A62Tt0cP5xYCxpSnVZojg9EP5jqxVI7BRb2pO75XqtCH6p4I3FzEU3vImjdZkjBkFj8HoB
5jx2dpO32XPF2QNzIrlmpiFYNwbSijENtI87BZCPKajm2KBfOZQIyZDCc9pjzFsemeXX4N0Xa9op
ynqMP8HklD1of8PLfZUXvHoCG56RusbUU64tt7wAv3SmMr67OGwT/MBT+xOkeIzPwuBdLVqXl5BX
exSKoVJ6uiMHO0coFMAjDwppiNHL7yZ9njJ2gi24LIJQToUgVly3TLkKNnINFFw4s6mGWpgtL2iE
4WPblwdj6IAWu7OZyZ3GWRH5QX8ArRwYWhRbdcvRRbQ5rLJlOESbf4JjqCF0S/1wX/z/X5lKsLV6
Gi7hw2vgpveTkMN13ckWbv34ZQZU7F+YIUeaRK8bRMn1ydoawC4WkGXQawsLSDxlHAyGvnp8l1ym
xPmBnhn0czxJp+TmpkF2BUxCbwuUSPJJhDsMGGONNWuu5PCiKs/iUobuaCUBhhIlULuc2lccuPV/
7yXhdWt5XZoZ/Fck9jUD30gWznEAdAUYr90xXnEsdUvWvysF6qsX9Umac9uOcnEiCGfB6cPPqBb1
pXOL8YtgbOTXFzbQW0VyIh4XzaeirUufPyANkqrgGaVUbuNfkr67JxAkKNpcrKOt8uiaalqhAaMu
VfFBe/4gebBe1gnr1Cy9Xlk4Q88/GhFC5b8dmWOhd7DSxSEnXST7BSi8J/ZVkgsdmnAcA10uwsFb
zBbRmvhK8risrzynhoqCmvIDx2M2MQjsB6hAwSIGIgxAPsgOzbzPolmLSANgvCd+GkVU3ZH9yIeM
ENcpHwqnE3D7+xlwvANAAaxeC4HlIf9NfBe5Crv5/wPKjJ6nUPxWMq3r7JMADhvMjUYEdmqZ2uUs
d/6vedZRmg5CVklTXlhwhTdHkCa1vVsKd4s6RohIGaaU46F9h1KxHftRXcNdw41wABqKq7DX0UJm
Kggyi/aTJcrh21vpwbv5S9r3dFGJsRrDnHdS+T0GhZnyR+JW7nCjRaXozORkkiSv/Bv6wUHXCl40
9PCLEW8Hm/emmqldIyYGUVeCGE/8G5ypEbUJEWQiEdokiPYEePW76A0GGe3gCcdF0BmYD3rRysVO
F+o/79NkULyIQTAMCGj7d16Um0FtFvrfBmqBfvs1kyBvRRMZRRndpMLq6QP5NFqakH4dbZ9q//Rx
92GDvZdsdxzRii2Xhismx5ytkOToH/tubwDwGWnNpEFSD69oGNKXJ0MdhnDY2iYNPZy4Jy+L7ddw
DaE3SK8ZdphdQZYO3iJ4wT1Dep1NXC8CuHkZHhsmeeC0ql214OE7Wi9uI3b2Jyrf0eAJxt0O4CAS
jBCsBMbuwpnzZ+AvWFQSq3n0+YxhXRim28Jl5Do9R8CXjQN/4KLagnZtyZvm/SMpYh9QSCTpoLYq
dZYQJQ/bh7Hx14U/q0HHGYLNbKhFeHumFByV4Pl8cOZC8bJN+pemx23CoZksOUWLIu/+UGMko/7E
LWJU2MFjAzQqXGH81Bm/UsDDwfIFZtc2rsZiIhHjNd6KAWdzIh9uHQPn8IfQTiCD0Alwp1vWXTUb
OPxFhaJLY0Mt+Y1eTxfT3O5YtOfqhznDXrUA6DWJ+VYLnpZfYnGLj29ygZ6A4nbbI9qWRz5pMPh6
2Um1nw4c+A7YImJ0jryhEnVwkk5vPWoYc90yVpCIfzeQulYWfywEIsRLLph9C+9fkZxtXxMYqKEz
NjPg36fbeNgAi11ehEZ/7wiKeHxgEVXZK6Yjo5ksQKq8dvgeIxYETkAjoDU2ghzzn9rqcDqqpR/c
7KM8Z80WYhBY/vUAqR/S6+83TcQYLtF4w82UX+Qq3OOvUcS0b1WSG8LfX+//4sbWET+rhPPR7f/N
Kole/Yg7IptGqwOlmq3bU85R7nI4d0+iQz22bHsOh2Lsb4SM5VufFcO5HU6NoH+eZdmvyLdppVED
nqIwQc00hxQR0+sVAU3bT+/9N8THkQ3cFJFM63eXSjencuyV1Nb5W3/wTo2JG68UWuPQfnS91l0o
h9EImOZKWfodaYRkbwam+d2/nVh6XhzCF/BboDbrR+BefVBd9xs5Wp/Gz5OgmaoQAzgpUwqBspF7
PiqLi2sihsyrykKGa9YWIxv47m8D8DuKI/PTAFE6tPx8h5J7wiXyOKdX9XfR8guvsFFLsiitURMX
SVCHt0IP+5FR1fPAiwEkrx2bLgsWAPoIXAAOQF2ac7ZCy6WIQgPIrU1HFu8AuwcZmY135T4PH8mc
vJrUV4S1fut07hwtJXdghBa0oUx0vBzKfS32uBs5WDdnE74SERXVsfckxNlX/uthqhwr97LdkD9E
Irc8vJgZTzmvhXJ/2TZFqtM5YVxZyPLGEtjMKkEgr2J7+RldQVeV/gW7RSsAhvM1IebcY9v3X+PB
PE6D1h8Y+bR4J8qyZtGM3Nuvp0DQ1tjtnbl6o+GNr4jYhe/jKNmdhXmjP9dlE/XOm1OLlVYQlG8n
LfYQQgx+xFXnBBLn43lEM/TLB7OgsvwLevxGNaiIGfsVC9sl7BQIn3vPVlAzwoY7TfiN1N8byNJl
Vrh19RcBCiG4Uv+Kifq5Q8WH6bkxs5hIkihD5SESmyfFFbbV8eoZgv8xeM1VSA7Zhi1hMWCLN1p6
Uw87cE6cMyQgrQwjKXSachhuxUhkEX2BO+DCleVscCFK7SlzUHrfxHnDO96h9zcs/CIjafhsp1Kv
bjg3n5HuM48aavHSUzog5IC1udXhBwawVrR1/gS5r8twms5FRhbP0+Iw9vCY39xWt1KoxhFimkCn
uGmukKM/NC2h6rcEJvmDpr2a+8cQruB8fCqd2r2gn7vN1HLpRdy9ZqNkEk7uVKxPKuaUVAOXpIec
6qsJDWUIsJuFpnPLYxeK7cK+xrDGJZ7Z8tlK7TxFbdt0ir1X+c6g+ctYLG313xnxpy4RuyoMmVxk
15SgH8vZm4Rv8DGE4vV+jKna/qWeppdoI1Ch/nSEFnu7zFclXjO9lSl8tGwr4R37QwK1L69wFse+
/3vhRCoSdE+b02MW3dbtpXVytkiemCeb3A8lb+yj2heerheoiSN/KbaZEg4Z3w4AxU0cZLCRC0vE
mU8a4WvhoFHh9WnVnIQchh7tOt88xC0OlspFrIfv1kfMOW49XOiE9fRlccpkFz6Iy4BWKy0xBG7O
T4CbSveX3JijM0+FAQwPDJAkIg6y+ZpONOguE10m4mfVzgiJtMfXqCUox+OFKv2EV/EVDkC5CmCk
xxhaDnHMDKJ/a4JakVsNJOGxnoNeU/WuQUKIKYpYucxhprFzsP2JHMmV9xpS7PhshiTIoaPMYev1
ERTdVJfSF+OSdWpJeBYUnLmzZjTV4Vx/wN3OVjKiuCtyfts2FPn/6ZGUlDbk4EBSI4XfLWqTJIGH
YnFaEf1XK7MlJLTPrBw0pNCthqVbchAFYrYU8MJJLSnv5F//1u/Qj4BUvcOyTktNPN10C2oM6hXG
CWhIZ+D02kfTZ/p6mI60zAQ6EX/i8j01L0AjnkPOl9pzIRxtLpYEK3hCUQw48GUgBWPk2YGGLgoU
Yefk5cBByLcXMqx4qBDG4dEqAYGnKzyDALr70qvZfc33AbrtOu3jSPU81bhb9oSimxmZpt+lL2Jj
LCsAFifhcg9V9cTgWiz/hSazIT6BtGoorJlxp7TN4LqrVLiDwHVIxXVRduA5qWpsEhMbCm6d4UGb
vDuty2KgrH5HRD+KqDZIEvF4uCrhUap56F/96UsFnSoZ98HmH2BJit0M8QfOWpEXJ0IlNZPJ3t1O
eldcssv+15RiZCWcs+a9AIMZy8nTysVX6dssy69MCKWY4v8PamPUyPzXWUf/6VxHtuwv89WZJGna
6ivx3XyndhqiaCnWtdG+rjSmyJa1M5OKiNDN9Y37I1QhRfIR5BAgBDfHKVa152v9VDakjJ8jfLnK
vFVn32V03AbhF/08GoAu0y6l43+SylDJcoYISaqd0vEH/szxBNsxOZjlEUrT5I8ynxFePqA/SNxB
cqUfBRFfj3JAhn/judJZwGnSFP2Cs5WnztCMIfxOttKbIpUxc2+S3CTEpgm14TDLXZWfrcTEzwBm
JdSRGnnDhq6BSDQeTuDzJbaEJeA+GXwWU3EwUylHW+/MHGM1Zr2qu3L1K7Mgw1urY9DJnLiAr0Tl
6g4Nd1kTQkyX9gdVpqkcmDyZtKgKUSQh1N+hFYEhYHFG4KpvgBNznyhzr4zQG+nmh9iWkE3Wwrko
8UMK+vt3fcQEZsDm5C/RGxmP/hIanBXAf0SgNFNW7X6WAl0DQkdrE5l5WyhVu68ZfBlWBYF0uSf8
9dj3jku8j6cD1MnFpNsygQAgHMw8wJhjuoVPQIshxNUp5WmRNsK6lczvquffBpfkpm8AGvoYavT1
qw2/jlQvVMvwbrloaIgw+Szmv1g5SBu4oCYRPYUSw7kSaXC1bCY96efP1sLkCSLHls4u6DsmkOeY
dmNMV/iLdFwtcFB0TBLRIqg5fxKyKJtK2uLNmoTYPkbcHGBnHiSrzxQwMtWPhZBL9O3X995oQ9aI
qPFrCDc1P2wM0PLMpkospZu19uwO1WEFBi9QRc5HJDTEdmdJhw2abP4K+Eh0yosjdOcbL5HFXvyM
/OFsjXWremLuj+kDKvGbfWeVyuRBuZZmhm/6yUqkPKRcjNRtQLOE6FIFhP+Y+VqyiRTUIEpjnR3a
vqYvRrAw159r13rYsrZVwq1cwdQ0TKPSDCjKIXB+a/77BwcDMZsZC9b5zWdDPGrL4XhgSXU72iJI
NFaFqf78S3roOBa6xphMqmjcGVxPGmq7LnPkTKbkcgZxnEz26b/I/feRnkbHOWCZB8Ylqhb392JY
DmOYw6I6kK7+FvmeHpUJ3wqqigjx7GOg7G4Z7KU90gdiUQpYTCLXrOvovdJNsj92NMHelTOLyPpp
2QyWuShm3PbAvdOjDAtmkBGj0gC8Hx1xex0bYFOofeLAAdH7NT/K6eTq6QTfUVneMGdqu00J4MvI
1wn47tYalzkKMDpbs/Coht9LKi4rDBdfK+NU8ql7TJcR6AyoFya+dPzXqeq9BCRZZSUFZKS/GFwT
6uayOAmx214ENRAnNXXM0WNOvo5cDoWPop7irlbR4me0QstiuokEb46B4/TPf+ugTxDex5cD3JA3
W9pq+fClVuFaslJ6ysIVpFFdKmJU/Z5yKsbchTrNqWYmLaaG2fPhHja3ubHbbcm8vbFFwarQbq6c
cd6D7OiXbQJNK29hvKSTRiuXFC2BnSwwMTljtZSRAfJL5bJbfmF6uKbEDSssc3c8JzVVzAYqMF0/
o+ShGSo1ghJpLIrugcb0USzt8KuwejGJDUgkCMzLmmsPHx8/+rn7mY3QvSXaC5MVv8CaIdT4SsT2
j8iHDxC3scsCBdZf4t9iqqSpFyAu9L8Iw/CBE5SULsR/oXFJmuqlQFboY+7CZqiJJ6nht1trmcG8
NjKi7KRV1uLZDO6I2/ukhDzU38haE7v+LaH6XvNG1v7G6k+i11lwwsImHl4095U5F9sZD/hyI2Hb
vXLx0PN+a8qD52mjC2rgr+bsu9n7nn7X2l22aiARXEr+f45Xx9nvOyJKoxp+oPLQTPvWpnZNOfnU
zFuxq8lVDhPwvdl2XT0rp+WPqxiydHPj19tCxX8zCpwqLyACJRAafRDv0gsXV7S+naknviLbZ2ro
aUVgDZPKi3x5+zE99rKaBpyMgqde1SS7qfWGQzG9juRO06v3lc7XquMfQI2D8u/vRY3v+WJ4ZxG0
bxIMugUrC2dp/azBuske4+NSou9cHPaymENul2hSdWU3muavxvT6zxZqasToyTfSCyp7Sq6atNFL
cgmmEgvxHb4OWNvrv669963o8Srq658J6khDJeuoqZZkiOpk/dsTtggbamzxdke44IGij3tX1iJU
nKzkuOFcgjKlqOFYqFPygoft3VHr32klIILeT5RPHgZ47BQKufTgCnlPOtIg8d8Nq3LswJ3wEiTM
V0AnKfOgtQLTe70FtzcJW5QSM03CbCSgUb9zJgTECy7pX9zhTECdE2cKhiCObuV2pVKxj3p/rz5B
wdM4vRUQpqHtDaIBKEG9HOqNqGtpnLrFRd+dpvC0j1NlslWjlXGnNaOo9MdrdZQFoL5vcx5IMSN8
KYzzMkapCdqlYzHy4izc4ZBDGvOZSOEFbqX9S3Fd55o0Cpy4gWGNgh+rdN4CLsjGC8occ1addqbj
3wnAEu8zZ75WXeFVPHdPKLj+E9MrRaYQ4AQ/yG+y039TOexugsK94V/amsKJLzqNXimSi6PRacV5
/obQjRV8hXahfdc5bFL1i9t4g874MYJ0+j7uvxLM5bvY2LtwH/PkgWyldN/O8O6qphFjzFzc2e87
CLmzrv0oN0oNdPzedi2slIZOU8ttVvwln7tMVIwIbfQ+SOXqpW402Xxdeb0Kafla44eQTLrtScR9
Ji1dJyi4a/ln2ylmKaIro4vavlyAJfh+zX3G25fbFe7wc/v2KO8m7YL6/jtYUz1PPyh5q6dOHUQ4
fXt8AVgrLq9xy1erPZVK8ScPybCt/bpKtULzq7gnULqgVkKZArpo1TSw8/UiaT1HAfMy+Uj0yDtR
LzmWE2yyA6oLg6+gN1vXHQnRClQiCcZn39uNysVm43+mpNMAL1HsN11nfJHoqFTRyWL6ZpDjVNXg
2TtGqs9YaAePIol6hOJjV9EJ3ERscNfDLFUFBKNQd+LpYwdUbH8c+qBlHArbyE2OM6GZO+FlxwJ5
wNJ2Xogm1lph37fdAARJzQNJSp9uACuJsqnyk9dbX02/bgKOKnNq+ZzH5Jtmn5QtLbyU31kqBcDs
suKzscSrKynPvVrlvwZ+R9zLWWJExQ9hUVnU67kmCYVMkZWsTe37PysVU7udhV/8R5qAmCgbG8Ml
oG3vgQ+mHxA6f8oRyqjnczFk3K5n1dGtdSdXgcqPBi2u/J/4b7t9LWk1+0A+M4Rtv9cCu/aKzcoc
8L/ATyVD7n/oKRRQePRL1fmtuJLJ/D1lBHN/Xcaq768kXvBop2U68IrF1RryiA+ZjaquaBGV9KMm
mXJ+eqaq0P3JKsx++k2ULXu+A0D1EEBApJMyJsEg8F54Xyj0bClBL1gClB9QF73tYOSuQnG/WGrd
/KxKDPTpu3aWSfyH43JNEuPHsdFSDuRkWiG57uTce2g/nWVmk15qzjO0Tft+gRFkgVl3WZ9jblZI
KIXmIQ0z64jp4SuKr+4KtSEcuGEMwD0sRr88lMdgZmslqjvCJlg5aruX5c0Zwl/9W41cOn1Q8DQi
S6QjfnzrVVeixc4fFen4gHePmuzWe1evi6IOu9tz62vIwWc7MX9lN1fGwKI/fKkejm0iT8YoJVdM
sbN5dmiKwABwrUm5gU34BnqWZDMA132Fm6PnMDdzJvPqJ/ZP37frvnHRdd2twfSwBasc3OObHgnw
fe1D1thNkoDpnq6C76/rhYfeCYJJcaoLGTVa5m174EhEcQF0gJ5l5IzACC7YW7T7Qzc6SceXVtFL
6p7DKe3/+w77gwTFb/C/EEw7OhEYFM+XPiwocqASn1WNhOqsBlHb8MkJNGAX83pqcN4hhYZHAtbS
A3xqhjmK0Nbs90bxaG6ozkODe2dX5PterJ9L/8jMci0YFL2mA34XFEEIGzFiHfTWqGakPUz/cICe
xAcytGWyz1MBNNNHKV0m2wqjYLwE35zbLANlXxJuuhG6FYww77zc1DHL71BwvQwjp7VAM8La73pC
4IRSpjxC3ME9Ybq60A/jXF3chKYKoeXW53e6TSFwIm0H62Uv37JrdDku6h99A/5vdsQJzauHJN7p
0fL2lo+L5zuA3jAIiRJglldJo1ETSiuz/gAYkjkYPv4vLsA64J09E0UYAL01tXC3nW66gKFYkrDw
A3sOmbMfkOA+p09Aqxso/qjm+EqVEp1hgHSyVP2Y0Ghk9aeDE20DuhlRit+5Nuf7Zo5uPVzJIzgi
ryiZ8KtcadwvtPUjGZTN1OZHjptiTLVZ7ajFlY2eaDwjCm0QgHP6DkhxV6MHk3O66LEN60gYdcVg
kxu2WdPAgNKlJYzBXJczxQWgvHmCJV3Jvkoth6od/1qI7zC9HuQbiwfneZNmf6rFNH/yBy5SFen9
UGA5phZKSubMmO6pjh5pHez3pIjppfhOMDKs2IJ1efSvTQsULD78KTjkPTTkl3KUZNjnLstM5rWN
YH4Ve3dOsgHS1u5IryvGEircVage9BLhNGyuBUl45GH0D4XK698XKjFyzmvrg1qeg17jamFURoAg
HwpUVrHrTeiSvGlXtwBkp638k5p4ckL9l9Q7R/mMlvN0uBkWN6+INVy1KLlrKUXkTvTazK9AfS8c
TW1+H1VMtNxxI9/tFjxG7lfU9q8M1BhH5LA+ihxzpi5ceYZUaFYaK10YMuDM2nikNYmYNxvwwsMW
ZuNHO8yaQqeau6h6r15CyQ8YjxiXtifIusD/XrYL+dodNkWncmIDJwFOv/fqdBD96NJ06j5thn3L
lYMMXQTiVtsPPue8FbLk+Br5gtN4KLD+jWAuZeEVcMKV7q9/2zyYswt5SgKVM1yrlyyN36rueOOs
Z/fSh6T8g9oM6A9FYC7FTIBJ1VxVJQ5ulqKujtBfV8CIktRwWv/W9UV3CaQrVymDiUhgY6dpX/mE
ccE5teRwt2fVYJOEBB2DRVezrzKWSH6uPgggbgzU1KnF3wQem7+b7GsbUPmfPC51DGiJkO1j+WFP
WxLXRsuJCFS5eAavSrOi/CQTeoeXHVKXSVQHfmHM0ma3U3voLdGhy7Tgu6TowgqGS5YmBXw/W4aI
sORyFTW0RHxzLzAWZ9ESBp1Xv3q1qxxxsGJjBROryEvzfzMbUF/0EesXYiFY3pEL5sr7kcme+NGm
og0mvbSKyroIJTTNNhrgT6MV7yZyA7opUlbckWHUGp+wtUt89eNyYHAy+DoDJJBmPRGAA/woRkCh
uqvj4GmC8CwEKDVlg4Y9kPbyfKC2sss5LqVKH6cjGKulwjDktRviLzfFB0TAT7YZR/7+E38K772Y
bfqzAY4ej4jD9YwnexqwQrtD0ogz5BFx7W22J6aVa37bDS3d3C6/djpLL1wtswNVaEOcl6BBUJST
bPeLhhC9MwzeVnCn6DzK4QB5uNxs+bydDARr7JUgtQHu7wsuKdeShUYgh9eKwrB0hnMjeZbhsTpU
27ZYGE2DYNidkmejLkZvJs+cRWZHiotOKgai0UJ+4li78bcO1vx7cBcftKKBe0p/gn0iq6SKo/Mm
XY/q0uDCRetAhgf1lAqTpTEQy37SdPTbw2wgT7u3uSUZaDppuIw0Uq6QiBtBsZXok7obZnJEgbfY
JMqg/8cjb89IztOvhxcsSDC8l6jbPj2q1w571lBRn0YkAvWcqSX5NH1qy0ixuWflXEYZsuPvzmyG
KIJTShui2gshenHJm14tI9zm/PxDShuRc7dwvIIHCyUxiOIos4bBnb+RXbCB3oy3zJ0jV3zgGUJ9
JqHtG2vrDrBqnUcSUmTUDHwwuvNC5DN3us7vP0fRr0SZhtoB/oHDcXeaU/nZLPQX5POMQ6D4Rcti
gSh5MyFd1C04YmwplOEDR8g1pQUtjQUq93GVYJjjDXOWaj1pGPxnquf9FkN7feXZr7wm4CvPtdKh
iEoJh78U+RGlaaFgjU2mRf0TedrT1T4mO+cjU9z4zfVsQxqsiMTksHvsngD0NWx2lzVyJDqHoh8v
Mb642wQwQFoJjX8azBsykuMas29/wXZZPAToiud108maoRxrxb6B2v63j0q0KPg2j8FNnCqcwv1i
glC9nxtiIm2zWIgUg+DD6RfL2+Ytr2f/vlsaa05LYwb/prmg+1q67aNf2/qWd53kN5qldD4WDZVs
kA0em8MudB10Rf0KgDlCOKfAHefm10hUKHoAlvQAp7zGaYVjt+FM/enn/d3sM3Z4x2LQ6G7oLdE9
KB85FDExtTmc6VvhzNzlWuKdTs5dY98KEP5LX/twZs2kncI+nooGKhbU+3j44rVRgpJ7vk5TK6FN
eK/S2QoO598bHFpDKWDgiWPQOBRt7DDFjHSUCzOFCE8w9llXRm2KPlQxaAvShYykYfPjCNdQSAvj
OzrP/YBerTYDwwLwn8U80CtaIIXGgTwJgVa+kHZctyefohNZJ1fng0qBWEQEpPDA8eF7VOX2rqyN
dsZ3ISOru0yXZn8rkv6ECbWXXa7GrG2DwRstoU5Qu9dxMJhm1PpOoO2gAOe+gHSXqvV989zFd6KH
1Ti9iELZKXZGuF83r7NyQxfELK6dMyP8E7CSSP6kLIpXlpxj3s5FZktNKgy4Y7p+qyhcilJVRzAz
gMeN7isInKU+vI374GINliNOrKiMBZN09v+v0SPSBq48qRhulnUGIExGVjJtQswksUwyetOCZQS8
eTJlidNhg1Fsu5UqhMqkLpIEc2ko0Bxe0tn8H7oNxr8j7nmeNOQKCNY4mXVwwZPKZshUxxR+G0hi
DY/MFZmA19z9ZlCok4bJxJffeEK368k8f+uxdVFvPgo9BfqrUL+x98ky+larZRS0DUq4+Yv9lB2L
BeqUGSVYYe/lv0MOyAn+7EZwCQ82PD2QE4qUdHriZoTwtCGd13R7eLc2f40nm4L4fd7Bf+hDlIe/
xRTQ2YT8U45l0mYKMGVsie2PODHCiY3Ig776bW2dwCIwdk33R2KMiE3F0RTRtDDne0A/f5b4yOSU
q6LPThSR7Si39kr6/urbiJb3p24JdnSvxA3N9GQpzL5jS0byI88uFL0KzRzJAvBa8rFN/oovwBZC
I52txLTlq598HcU1/K1o5JUDhzlo7jfmh3LIXC5BPE5LYFWSplv03IF1IzZZykDR0gYym+OKww1Q
1DyBrjCLMC2C1rGRUdpvV6Lipy3HYwUySE58agecVDGb1FCYvSXbPvzCJgsJkxq6Ewv7+YoP5Rxo
xNPf7VGt6f/x2pZVtunAerSuLRFT4IZ0zlWMbDYnSzPw7vn0BSt29QVR9WOMrGKiU+RK4OwuBGAU
SozLABxNYDivcerfZU80mGgKJdqsCgvlADBWzDxyOW8Rs7kVRhnqagDTYmvAapHyPT8F9XACSVAp
uSFje1y3hmaM6sCDrANTyOGkm/NJDydo5KLWrzD+PH1BirTZKhagPp5AkqY2dsA5X8gtOwdyTVg0
DBzzUR7BwJnWl821J6rPAzxVitFSKodJPuEEzvsadXp3lTx6zcZZHF4TbK3BYej2Yih9O4kuIttp
le+lkgQhmZ2ZwO6AfyyyMcwB6aHHScjFLu+YkEJ+9TbqmNyxhJ1AsshAwp47Bbe9qg1cBPMpjWKs
2Enpb70fsL3XFFf8dsrgD8YvgOJ3AD5LaY3FWd5V/kZJMhluoBFr/bMZh2ea6OGxaus1yb5XxFjo
7nMfMHa0oLSC9S2BvRJ2DhQovY5IZB9v9x9S3EEcxHu4UWdS7t0W+XTw3AOSjOe2+iLrt1B17VVH
Uqs5GpqRiXGrorKJmnYC1sh8I5k304NxEBFSfej5nW+IRb3oj9e6/kCJa4rbktIkf1BZbMzqXy2e
o5/7rF0n1KELjk9n7kEIAZj02UoohYfTIUlEnXoX7vOApjKp5RJzrWixGUNCzdmgChJg6sMr5ghp
bO+OHHvGTke6Jn7dazjJKfKrMRk5VB1RHGQNECiClfmP9fPtIx14TS711JQjc5lTIal75SuHFss+
doItFnugxxztcAEPJCqY4PU0/WDE5TT5fxAMBC1D3Lv06FaANTI83bI6Zgr63fMoCYhLyttcbVVr
uurcsu3yb2qozlkf5aFrbQOCB1O91EhOxGXYZHcVJZrO1xg//4z+4ZKHq2qEZ84i5HmUj4wydFOj
s1WZ1CIQ1nhYQsV+iYqFC6TQGf1g6fwKDWHrV/Px9F7RMUh416GIww+ounCJtBGMLX6R2y2BHISB
/QP/kaqhnmnu4a+WVA9JclfggbWUWzdmzMJtxF7ExGNKg5Ceds1aU1SpRigNlUpeDSMV4dbNFtlO
7dfrrFCidD7qMd2rc327zRKYFIHc24lue7SB7D6dNQJldRhABEI89YdV9M9WzJKkKAwgX3T21Vez
BnW/Aqsa3IZ4qHqv67k3z70KOyuJrD2DsI1qcGPUNONwvudhqCQmrlZ4OSc3xzlCz8NaDyRdG58Z
RPIwSudXjf7+L9es1xFD11PW5EqWATExJKlAn1oCQG6qJUL7nntLbRLBF9etg5PGu5wxvSmcpxrq
7xW1eMwU692N57gqIUIdQ97MtDcgbrZTR9UQ7TiHVJJLCW88VdeKtFr9MdKW40ekG0oI3ryJ8Nzz
1bp4VajYQ8UXhhfFedMXUURiDxFFqWU8gc40bgP/a7ZgvfegRB4d9doarTGh4BVmCWgQ7Th8zAMq
8MvIf7Jm8yge3qoW+dAVNtumjtGQ5/u4UGPm10vEMWAjguHU4J4RODc8Dypl/MeB6XNCci/zBbJJ
HDUsVfFly8uVQNJfu3ehaJ0hzaBTz0pJYroGdXlsW01N05UIlKpmFISGukLl89zg498uiMY2Ky9K
axTGPhCvSx7Od20IXKa5ccPqAyledo5sDaHeIQbyydCT8xtCv6L3ro1gVt+cC7+PSI+X1k2B0tPR
BrDW9fFkWSBq3oR82ebTMgtEd7ithTFz5zjKEXkkqELw+WWyKoQtPyO0Vxv+WbifCmc2MPJdMvtT
b/fy/qA7NUElfruRvaxjQ0E9QH5BQnxMJIX75t+M4l6kjKlEMUnIcbJXCSYo5ROD6t+bgfzk+aAp
PNzVvJcj/45F4d4yejM4v8Qvj78ThjlKjFqLgV7B+psHw0oUPINGqhwM4g9EpaZIKr8djNs6WC7e
Q9utEQHH+sX2GNgMl/7l2PQ8f9+YInOUx3NkLcoUu00neSjB9CN0x0vjneuwpU/657+lLVKAXjUw
t3cOtbigCcPiuzueZpHbrZb4d/H/lJ2gZNHAL1uB79ztdi/wW2TVsZbPW8/mtFB41c5EeRIkhcwU
xhiCjq/PQLiBhCd8SYNQ0U1U2umzJc/U1imApqYsfFy0hdIcgapAX09U45tvpwl+CS4+bL44FUbz
HuWzqcOu4lUA0SYtYT42AmhW9TPSda7wrFgb5JqbpD0utcOmMM0w7z491goku2iP6sqV1JkgAIux
AgsLDokgMsVwKPo+jhkktf7njEOcjLmDvq5qZe6kMPtaPjE/nVYY4ROJjhKX1fIQsz+JSRbz2jz8
72pzPy729ntsw0tljkF5SRN5k5hxmq1i6IaJH3vBC4BazGVaznzsbRV0jYYokxHGn+sk1x2fLvlk
U3yHUbI25n2JT3J6mgfwdBcjuluJe3kLVpxHQDCw0PtD7MMBgHlHrvPisX33Mma2GDRAo754NvOw
0SnP60+VpJdPu7Xm7Twt09+YZ5/hS59t15wr2dV85D5Of0R1YZW57hFZ9UMFCrBnptjhnvRQfenH
HbMIitcLNOsG4ZeVNPAXl0lo28xUDeZt1867hy68NJxQWJ7EFxzutI7I4vLfws4+u+8NdnsKy+AX
Ho+ZJvAZ5vpXsreCv1SD+wg2K0P1bcUnhzIHZ4meUw4+uJqRaOIrJOa6U77vFo33gQE0LgE9S3R5
ixZDAVxNThhO1aNMgTy06swxgiJQ2UMnokME1Jk65bjxH7DqbEs7KmsQEl4wofdG3L2z3i9M36n3
4E2C6WAwlA0XNiT+eFR51zg5DU0CnbXZf+MesAZnxq0OqY3H0D/9WyiLlWj1fKY708ix/viEDolk
HbTu7UGZPqFQ+bCsLTVhENGAYykdlqY2kCizgI5VV7ehBzCnr120W5hrYIXV5ZNGxv60rv3ri+2M
2GmKusKPCJbBOHHFKhYkIIahSMD7zjM8HO3Vou5ukldm77rslck5ihQs88of7d6ceOV69Nas4qRx
cN6gt5W38+Dqbp8s6BjNrrSsPFW2OBRzt6n5Qg1WAAshP7lddXOCdGGIpBtL7O5Ta5YH2aVi130o
WfSkFyMghn2bj8cMg8Ku5Yse4MFH+lKGUj/uAZwKVxe9vBWoxh/og5KlXS3LMFNQMS2fltF93QU6
L4HUsMoO+y6+rPZkr9EXaeP3yTYaNMUuHsLPAIm/AQDMNl0fJD5pE8cWjm0JZ7rbVTPpOAB+5yxy
YUHziAiAdM0Cce/xBdgNJGiITj3iwRXaIjO+JEQov3mB792QIua1qp0NO9JCxNyqTbnOoquRpFbc
aC4Iecx4vAWRwGvj3jlG6g30DKnkFT3hTUU49TMPoWGBY275DVJwpYRlKGGtK1mZRgy00Nb3H6VM
bw/jiOz88ruVGA5ohXGOqtmsTYmaOQOf5WOUvXfRn0xLtxbLm9QRlElHLBsyW/w0dV+w150A1Myx
ug68bAJhl6bbhaLWxB5g18iyo8X0KT1sehkI3Jsu4ciKqzdzIz3jFqtcRF5jFvzldyzowFmR0EI9
6R6z+MDIzil+tO8z3oSApPdwJE4e8JgW4VrZutCIcZiAPzwLx8bP1p0MTtiszILQ9QjQLqmLsJVw
me5aa0t5CuosRz7cYTv2i2AfjwpIsxMO2aVkhlCKXIuB9kFkupFQl2vCAUtK/JqiPzwAk/cIuZI3
AE8Y0+2+GciZuQh33ZlLFrJ/qmMA42gNg4FgBnXp8HdDYxdKJtichZF2nAz4lFR+RzyqLBz5hUI8
jMKN1+3Swx68CweMFAUWYcD5nUSuNTzQdkOdQ3sQ/8V3n5QbAgsRL4qv+K3Ihv3IWHnFEgKRSmaJ
TJBYSVK3kqyQo3K82Y09HCxsiYyYCDuhSILFV4wfqecLzsQTZKHDiW6OfeSWNjVgL0bqvOBOx0Kt
C1nSongcvEhHpT3d+iczne/Qhp1Ff2AgK2EBI0X1RMdhXZO6YPACh9elP27XDIUU/pQ81pM04T3l
rEwpWUxqGyy0Maw53Ob2tn3g3zqOPEEOdwEOJQDISXL9rJwUbuM+OkT+CHm55XHYMsbH7UcePQMt
tYcJj2ouS+wy7dT3twqh8ODQ6OlAac2EMBrnO/JOdkBdKQmMBOulNQYK5Ia9XxXjLXwrTqeK1eFy
BwAC88wjQxjX2Owswfl5yhspu3TCR83BRAtArb7HGZg7rG/jLWhtD0/NncY0kWRxEZaMGsRGuwyE
+oLN5E46rahPXYIApVioBMrRWqzW5RS4XE89QxPuc5lR/DPZ/KQqotgAZ3KXm3RTgshe8/Yp/jR4
zX+CshQu3MAVYj3H53mcHWgXbQb7H3p5YCA0TV7La0hK5fs8DHo95n5dIwjMK8sDwO6pBvNYpWu9
qmJO90YiTxYcjasgujd6NqJkjUEoemMAQnqMBeNC66GLg3X4ipkfe6Kl/dHx9laP0c180bGQd7z6
yh3uP5Uz/h8DvNxrSjoGdIlMKrF4E2weTZ0uuFvqzDXL5Pimw8oblPpV4Y3lDvOl0lyuQgB5O1tE
xYOMhcpbMt2wmR5ZmlwZYTtYavmQ5NtXHN8jy+Gchzc8sEeTaedBDECAGo6PHNl1tKe9nuW4m3a5
Qv8um/dm4HYOvMmqglkJ7J1Ye8BMeaT1wKeXvzqE+aFJ9cp3Rd4PwBWMPCgBnKV+DQ1SR29sCpxm
aUmYrhus08MEW5GcmbUcV17uOie3DSSMCbS4YCTvKZw/hhzD29To0T/tdZ115JHBqzEsA1CGJ8sc
BA1e21fMCUAthSq7c5iwVvnt3pL3MIupcDikRRmiXo7AFfmzZuH/NXljiHdyw3haYvKGBmkxXa30
E9ZfcLQyOr06uH0geDhNaj9273MgsLXVgiWd6N/eM4Z+gSmkresxGalsutsP8M0KnGTMPZhgQJd0
J0C8OFMPayeJp7v98djnsud71+p8Mp3DnGO+JVpdL8vX+IAsrNeLHF9g3iEIjsYlGkNxdfqZzoLj
XnwYVXX29VsEJHUzuGOQVRb055Nu73DVu569E8oSvRLTgmkvCE5vcuVTnNue/xOb/umvKxdslHG1
h9fWqIiKMGq5oGs30fVNoBAEmlCR34SYTUsG8xcyre2B1f2qZZoT9WOsJCs43c3WPs7FSwsCuoxp
fLY3QHfvI/W7xahqvUaCsQ8iojlYXPPCwenPIbIVm34SFR1hu2WJEvKm6Zv0JXjxicuqH5dHiDS2
4GZJoxvphgkAPr8kniEW0GBcBE4hAbxTe+bdSqfyR+W7qzVlpMFAvTP3xl8bwePp9mDVVeUnT4dZ
LE4IhN9UFKLFcfAOQoGOuQUN/hT9IJtoYO9c/EHRRbpsNP7j453T98IofBk7n4cysxPeDniEyPsC
pD4l53CEL0F5wYTLyZMXc+cESRTbbBqE/ObRomBJfvnqswIIzDoc1nc5Cd43FaaGzksqM37ovuzW
J1TByhMDeVzNxsZh/ohvGw6YbRlHjkJsc70ygQzZtDEcfoGFVSJFyyvh2pNiQ8gnqsgFjIAFdrMt
u+nypNMHiA3Fq89OYcnFNtkmFZ3K443ohO55NF3+W/HSpQjRxSVCWinI/RsO+4yjGUujaIZFAkxG
tU5err+HM5vsvyUqOWBdWmv2IVg8xYbeo7gq6yEriLcNWHHphjxFnGEox6wiOJ4RpuKi6hy2T/+x
cl4d9JOLkZmKDVl1G2MV/NTW641JxKRS4Pou7GsGodE3P5NtOLzOLSrnuqYALsbX0KSqhh2nU1kU
bzGWU6ZZSGp2K/+OgY9zip3RlbCN/rGVI6dsZ5AEQygbRqmXctYsoBbMukyT6ylMfZ60m/5WyUnv
AaSVLoy7DwZSDM98mF8gRmsveoCL/XzBt6ThQckPmWwaQ9I9rNAbEhhAtN+b9Q4kRqYrlwohTnhV
kC1Sa/mb0vEqsmTK5Kcakqm/x/OlsBreAHHdozebwylTnlICTQ4PV5bZqW8n5MfGq6Eu9G41sZqL
AzqZQ3tqROmkr31e+4+fWNz6R1wIY+Fw2j1HflqVvjifwvgbq63j9TXCuUmKKM7wpenNusjG4fyK
1gR9QF/JM9o6ceIfhUI6tlg7bFXzwHF4s5Fx7GxqMk6Lnc+LWE3W2DOVBipCWNKtisZfu1wIBK5O
mbl0EEdqdIDENg5dO9yGg1JHuVudT/gufAuLeeKVbmeA4js3e3BBzhnDUt7neVW9n4BJAcejyjAO
dMI5dgIl9e5/mLPDDcUaF9X/bZU5m1EtTdDbWaumZn4y9RKWYgVWqePn1qSElnr6q7cbpMWDEnF0
liHFPYfmErdywhH3tMqwbh0s2N+FXXjUXvA5IMhH2gN5uEd7JTjsv1qLFFuSImybGbe6bZVNH948
S+Ur/6vj9zD4oSbcae6IZSHoiK4dbIBpXqBN5oTg/7HhMoZAZR9OKyM6XV3HpUlxyZJdhQ2VP/QU
NUPLwwaQMyzsAQMXcbsyvvPmJ1ozz0J0UUD0VwelPA+mC+KEBZXRGklf7T8liQOUVa+mt6ZqgGH9
FSb6Pnslu95PDyor2ghJ/g1em2ABrc0s2GGUsZ1FgeY5RoBpqBgXm1ljDA6Cx5byhLum8DzGkks8
CGKOLUZwPeG9xytnJDKir6VWriMzi+sEo3F5bG8Js3zDluFBexhjvRHRgLl3iBQakh2pAU2FqVXx
UyNI2weY15CGbj2Yenv8Kz3clU7JVKl1AdpUyUamHMR4zm6TzL295ozA3RvEKyDxuG0PL1ak0jTE
DQ8l74xtbZcjhd5G27zFMabZeieXYeUF0cEntR/D8bP6BA+Or8yC3m6IRLS6M9dHkEl8bdKICVUg
gcptsbuEGQh5+LchqmziicV83P54N2TvolcNoLUfPdKNCCN/xMx8oF0RP3gEu55AGRvAIDuQEFKu
bWx1rTHMYFZusA32GJosN3xcz38/ODKjj35QmY1Sya/wdcTIgnFexg7VVK5GjqSEsRSlKjXqpG1V
lT2AtTNboZs7imadaO92Z/c7/vnLGtT4HcoJ4dbNxR+wYrAJDnSInIoBZ4unUrF6wMiJE+aFaTi1
XQwVQPdsLihE+7khXM7wEk3NIZRVLiymdpqFVzK3F0uNU47bHr/z5bxMppxs18nUT8MMsR4KWNan
Oz58RHGnqVpLzwjjfVJ9BNLpBueKC9+nn/KSFzlOT7FJ+4Fh5l8EuZ0GUrvpyjX42kpV2WkB4fZl
1ZpZIlmbUFqsOYaa7IR7+4d10kxSi8xtqRMZVN6A7I7YdbjDqX8n2tX8siyi6l9HRPKs0dD2Z1Sz
WJeZyyuwhG1JbnXpSmHDr8IUaFl1IxJFWJogh4WHh0RJAiZI5mU9B/IGI1Wk4JRS/Xj5x6kGMm00
ijXzcpPKzOzSMr7hLRQnAaF/8w243rdEWf7fO8YK/0VKm1cOrcdBVj0LLxj7vbRj09rRcV6Gz/8J
5Z669R2JBn4Kr3hoUyB3fNZ4V6rHjK53HXSmMyx535tI/+nreIQHzrwLC4UfjXBr/a/rDdME9l3c
okujCJ+tHXOjTnMkaWpoF0pXYHe24hbKkCiZi3jA61g3+XpGqGZ819KpiIMz2VHkVJC389Q1fAao
g8jlSyRZXLW/wR7BR/LwMOhd4/OVNVhtAXpARVrfEvdpbJWhDO4MLAej9ry5CSWUJW0NXpNDwWbR
Xvj80tgvXQ1gzhR3I/7fcp01pkUtHcl9+bDGgy5Qfv4cvc1oSY5XuReLg+MmBbAeC6TP1j8Rn4GW
50oJnvsUFM8uxmfPuyjvzHvl+02xNU7uRH7Rq4dYwVumzftyVpQSzQOuE9x+LUzEwtCn6fdht17I
cCSCWB66XPDQ+NGnaMGTYXUCb6TUldmEMQe09DpDY9stlmGDlnQ2/IGZImVPG9F7N4UPOIeaQZm9
c6ztG1TejZJZGMbyDdzGj4klMgIVg1BJXb784H4IgOQ4WVuyNEUYALIF5S2eoRbjXaFrZw6TPJc1
DhRXC+/l7S3dIMBlmt6gfOKZzoh9oZnWYS55n85kuTJu5R6uOHKoVJHUJUnKXG4e5I2a+SeKwURY
bSk8Ljs1wuDkA0N9KAh0Tknb83h8PbZxTHwStAalaXb2tzLo7KBz4k+o34VoCav2ENo0lHT3VQBP
Dl+MvrBKkGPPySk35CbSrc1tASupTJQUrA7uqPPpxMg2Mwa8bfd+mBZIGUIj4sHlbD9waX2qcyp/
0SvEwtWzRB8m2w/ps3x0W3ljl7TiwL/kDF6IsepxgYWuVIIUfA9yleryovOvUBR4y1Uysc4sl3ac
Ws6MC7qGB+ceWiWU/uTsvOoNAOeXwSJ9061hoXpXTaEzskgJoz0P86FWa8kCpH9YRQs/MT+ViNPj
0hJf1ulAmU1t8EqiV3sVTbAvLNlIzO2L7/tUKgngmxnlsmkZ18SmAuyriceh4+K5/QVhvf+YvjGO
7rwavY3qlQx1HMjLUc0wvUucy1+qypGkrj5UpxJSEuZ1E3I4u+eLQHtLkhqzZRudpBB7B2ghLZs4
LkrDrbSQtbTitklaKFcY7yUOUDELGPOADOtjwI3un0FUbCTlOkJMLEn/biQL81Gejhwrn7n8dxB5
sr5akLqtTduIIQlEMlGmSIyRcN0jN3w51CZbXw81yfpzjdru9uydlhkuM2585V5YnAbW7CXHDddr
lRW8Ko71Zb69CKziwekMoiBOO6LkpHzDyEtAZSX+wdYyOErY59BCG7YWimCRPCMkrGmt6ycmMCQZ
wQSTUPZ3qbSg+C/ySJU8tyuwknSWKs4B1ZCWTeGmzTArmS+lTUKBeEoWvnv1ywzrzbEl6Gj2Sd5H
uVFNg/svResWC2yhnaBRuXdO5VnED6ubnaEqmZYw1X2X5+0jHRwlgLeAjYNE7BcD98wEC9f8HCe+
3qTsBeoV38t4g+JMlNqE5OpIKLeO/IHRsgJbBUKRomZjoCE04a0YG7nAUQ2F7fkR9Yf9YmrQ4Kk1
tMvfSAggllh4D9t80fFuMA0TGerl4vBO/KOVHlC7yHFJdYgEasyXFixkPrSM4BkUJeEWPLp6a7FK
RRfG46YdPumGGZ5q+xDZTBz0mZvRqglWNp0iXqLfgnwigTskNNejaJQxKWrJBlnwgjSdRv9FAO35
YMfom+FWEzlY/TVwnJ9UKpyQlUgXlnPXm+1dT8ZgFmPeX7s8FTETkFQmcvhmM0w92GwPoL9qJwd4
FzTFTNtkh3vmf0HOedRWZNj0elijdoGwfPEJ6Ov7SaBADAIWwpe91FHYl2e2E+gi2HZFuT9JqcES
Ll2DmHrQsliU0bsmRn7dLq/4e5dmTk8NDy/Fe7FT8rNVIxu5b2ByB/N5A5WCH5sV3lwcQhxKkrLw
+Y7RQJ68wF05Olb3qIHSQBWEmI23QJLl26Cxy4VaTzeUhmDLZ+ujcWgAFthO/lcgzyvzuQ+xpgQ4
N+oIz13WAV6mwiviiyAYWuy1UaGzzrUsEuiCTF/uC4N9IZmOGIkd0Z7ZoVWRJHoZzgAD7viv8+DV
0GtVQRZ/drqIWYQNt1GlOk2RnzGYyaWzlKQNpPPr5opyHEkOin463LF/1aXWGT2gwibwwreINKuw
ZsZlC8W+oYcRxCfktfR718mAsOv8Z4bsGUBUD7+UYVItj1O609gxhjDHZ2JUx+2QUgXH/AO7JHan
iEdwnLiiFpAsAWAGUW2bEALzcNFISpGLJ62IwWeBhGD4z6LPxY7TI0vVsdxg/bTATs26UzBdmv4x
wgkB3shpmDvMVwN3RXtMxgPeaiAJekJnAF+SJKYzaao4KtwPWVH+ICNqH838DNEhgS5hyB7vE/qp
8ygOSRDA7YquYAjFp/IKD0ADNw0qImytQti7xNG+GBIfkuiMlqxiFoajCYItduKjxkS6PNIB//1Z
EWAVy2ShB4z77/U3nzKUGFUSGQQ5tKe8cno8+lwyacpXOnT/2j2yf+zHkzv0GhAjifu2Qzyz9inj
VaFApYna0uGFLIl281p9EOqktu6wOoXrMv9ecHPSOhgJd0W9njBL4UW5tmnPwaI9C/4K+Hi7A3Gu
uo6iN5OFL5goRG8WR1aWw8zP1sRif1z9ETTuwfMBTaelKeMR8mCyxfDmoqTQwv73M5o9WbV32D5R
URV+UyHIuAgCD2lCG1v/02p0pcVwtUIFy/r50bjbk56fmiKF7CKLh4ZkvsI8nEi1wmfFUhi0Jh5Y
uiOgunjdSuLqocG91d2UQoy/aKtqoZj9ibrhhBi8dSd5LCvu327aLibFiri10ShG1dIl/Fz2CEkp
57KnDTyQ+rUJ1p79FRV5WyLXQadskHbgy1wNQSHdx1Nzo725/yPOlkVZ/L/EW5mj2Jw5enAaQ/dT
AGto1bfdIs/veYIWjACnmKqeCg4R0kOtSYAYEE6pT3fubz5iKmzRqUSXGEtzv7e35/JVDo/PMo3I
uJK+tarJm/k9OBC48hnyahzfdpJeL/JwsSfXZM4CpFS3v1m+LAzTHb8Lz/1ao0a+gGOKSzYMJedC
j8u5+UFKPLTszP71NcOPYcDUwyQgCEhUyHXwnD4ug9iNAJO3cDnNGNphonrjonmUySg/D1fsXJJB
08PhqNIhXjM31xvRT1KR+47O+CyDacQ/nGxPKCr9AXygPdZdFTM2zCQF0kxGO3IwsZWItkeGOMBX
FJxdRgaDGmzdngSu2SP9Uan8hOiaDyg95Z9A4zzSodwCQioKr4PBgOgwS3rXqhWshFHeW4lWbF8g
HcMxQcifICt8qvfZy5uG8QhrHuEhRxFmgeSbftm9HTnR5EQH4vSIBasT1FauXY1dqm3WUrXS4Y/r
YBXRtq+b9pgpvlXxcjqToCDA/SBHff/6x7WcdXHOrU++g++70Qe6QC+/W0L+0HuzydaaixipoKHx
mk+W9SEsA7OIQgjSAvLC0oBXllDtlNAgZIoUJ8xth38CV1F4r6QPdnLL1ybYk80/tN8MWuZjOPMV
SIqYB7IEJmaAiBgV5QV5g1iXZPKstXbPt+V68tL+oGF5t3ryUOLV56UjPRZ3dzGYYexjLvjRv6nM
vOokQgQ9S8HVG4GVlAgVPlp9AfYwcw2q8ve+9IVawLvMWr0bSuz414etNw4R/yf6j5EH6Ahi7qIP
FcsuSn2ajSnDSf1iu+/S2D/kmJ667XTZ+JvneklvgVgYnsS9cDOS2onUNP4mMWtkVORAGdGvt+zR
VNEh0Msbzg89yc+KL3CJynsj8s34aMqA0aWfVmJL30rFQGDTzYKsxacx6P+yQsv6EhphQqTBPj9Q
4Opb1cl2sei8QTLgmxogVZa+Us14s4cFJWn49mgSi/Z4g4ORO4bq+AL679Fx+VqDDQIZLIaoCzcP
zSu2BPIOq1h138QSENZhBgyqRmXSLJqScfbPJm3jhBPaiib8TR8tCbBsl2/qvUGTS2GTcqHVGonV
YE/IFJoJ9m1kElBioROq3pGZNArCOLWdoo3lOTVzzkgLIj/Pc1CQDeY4u4vkPywCJGr+Z4Jufyt1
zIYaoGhH+vPR2beutHL3dHv8U2G8DddkGhvwx1+ZbzjyyXXaHXBG7e1Ch6NmT9sbaKzM17hYD1BO
JCNSCCg4JYWhtrQdXS0gXyw+noPX+Py+fk7SRRKEindfzJgTOUWIB4KzLXw9NsJJfhRwXj/xUH/B
oiQfvf4UZorxpPrQ4960WWI01QhkrGppNmCFSIeQin2Lyu3a8ZDahTfuhnaFSt+LqtMJOGWxb5Ew
qmKME7evrB5mglWEK26dPn6SeCHo+KjkEwR/azbWA9yHKZgJmm9htHOQ1ZFH7jowAcyCW2kqB3ef
yK/Q+sJGDf6iFm471nbysWjK/PDJ0C1sYy0fKdAjmvvVyfEbSrUTI/Yg4GTyG6KQGz3oxrYb5LC/
Z1Ol6SEHBH6zDeN5beTb20w5NH5drzzpDjdl4QgrSv77kpkFcdtSFEEAAvI8AYc3ENQOj05fGUr0
zSE7xNHfvue+XtYoZQfhYuvg4EYoKr8krFC0Cg4IwHPTAcvdmWu6BCkRVaiRxS/HsQRp5JnGbd4h
TM9hvPFfIFNOloH+5yoxaK9g3OdggZX+uk1yKJiq18KpE3HwN0DhCJaiJ+r+UqGDFfjbjP6GwKJE
/jAMro68AXdnGpW7Cp6WREL9uZHltO88F2Vk/WYH8f21fboe+eWnOg0Em03kH5hTsRjb3T3EWMxn
988+Al1GGnibus2Ak0GQqDbKxOHzpg0a9oclPCXI3RK69tAPmJ0foXY3c6JLT5flEG3K9gVUkNbc
OnSDDu4ixXKuoZtju+LUrl6s8U5LNr+KIoC8LqfEhGhF7MWaUUqYrIskZg0xOoJekL4JA0KBVdgz
imkSXB+4QnLLcwOttNQVSWbjDhVXuU1OTpvRymYFtrXlw9DUIrJBaZvxH0WcNJFWbzpWk7rCOs3c
AMJrCOoESsHBs/18Z32Y0Sz9OER14TSp3zfpNPkAqs8r1lULrsBLfuTASx2btkZLl/nOApeJUWPk
lKSSXpQCSuz5L2w20dH6mMilJzShy4NhCPxVcpW/1mGUeBiEbcd0lU68Sf2e63WkNIWI2Qff8xsH
V3E4FRpzjaCLif3cKIJIVGWIjFrXo1lbXRk2JIidDBhC9nF6QVD+ZH3uULiNXQL9Ylfpnycnm625
nZciiJ5pFhnppanl4kt8TQ+og5B5xPZLX/UfyiJZoDLdi8Jj3k7r30p03S4gqUqbyLKhVU064c0C
Msds1BOvO/N+f64kGXMQHh4AbRHbzV8f9F3GcRXEUWa0e7D8slE/Ye51vjBVbvxu0LBc79K6vcCk
Mek+XR4NqM9Nce1wI62X+5/9Wz82tLaY6tnx2Lwm0vls42wqnwVcdpbRUNvsmq0hcgKvOtegAPtH
2obLQdpZHwwMI7vkZBqP3kV3LdXaZP0lU0jlQpsImXlM9HMr+q71nvRba1emBI1nx0dWkoidDhnQ
A95Sr9ZT1b2kILBclob04AigQbaZpcziK95GfkIH9RURZjkTAm060vgJgLdgiIGDcG7Nt6w3wbID
I/vmFlGVs0BTR/wszI36vuBcYAUPUHOelUjpuMELBLHjp/kv3Wahbl8cTqORvFx+IkiPET4TmGGT
P1m2Vggf1n9+A/vEJNbybYqPsPJcQOY+bfs0FC0QBzJfGV7b6p3ZmNJlNIUlwPIFMx4mXZdqCPxB
t89uimLQ2qJeg67bxppKv28Ov+WMWgI3DIrgCjgEZTsdIHucQuonWGzLshKWo8qYEYsVvkKVJYmd
9NOgqIxBXMQFzngi6VftrM+2x+2TJMgwQcc5hNpViUCU7ROAA0wdnqyGhyV11xeWDwid6dA4774+
1txSMboWLxj1tTOCpSPhngMOPx2R5BhJaZ2TGKxWOZE52VohRZbmbzdc+oB9bpdjLhWVkDJNktPh
L+HdQ9uyRSlizzIicT916RqZzPXRaJzczzfkNC8Ziowf2KX7iZqKXau1yvTnH/0xVe1aOCstJ3Hy
Cv3yztVP68HEH/s1kDGVHOh84AJm/gwQGijz8n2FrcmmQdCat+hQ9hWZEWJzIVayZaLi4/9DqyAw
0SXgPmgstFfJB/BhLOOxjsOaWCXghwR94OHaMEgStwlB0DIeorQ8edTaxD5XZZs5La4wKK4tae31
TsgHKCp/dd3PsSnpB9gSRveB8CifNkyVZsFA+Alnd0iUUlKEifwOjFtDVMohyO4KVnHJre1Mu4rt
3JHLoG3PtCQxbwBm6YS3voDVgN52adLR47hrHvaOrIrZ+FwaPYp2SOMGxEmbEGiWWEXS50sZNvma
RQq7yzwEFLn7ESmVaiXgoNCnAlfnzdsJCDFtU+aCzLg7VRXN2NwgFtNdY3SfNFsbtfanwcSpKUmv
J2ai01Zd8vKvmSdMSGNZBCTrExegKIdlXGm5yf/yK264Z7NzGsD3+eddKCAhCeEQxKx2apF/Gt2C
loZ95D954/Mo5tgvyqWY1CkqodbpIYWa8DXjKIWgzghmfQTxNusbyiofw1Ne7vhCXoZTsrVCDffB
m7McyoM+JDeI8dpwNrIexPRHXmaRz+JdP4A9eNrFmUqRizRC32bRuLMoWo7rfwG7Cbsc/wqyDWZY
Ix9jp2eb3bIJalzkQN8yRx26G5cAqjlF+Ag8se9ybyk2D8/qmiAV238SRGkslNFsjD4c4OIX1d+F
WOy0QnJn/Ng7LuzIh/ln35twyifpBAEqxeku2Dauw6lbSCMRXKOwTS3rMFqt8Vp63Lu31B+rQd2T
/Iegaf1Ez9vc+lhAy7t1e2Phm+d79vItCC9+WVE7O+zK1kOKEg2skNtZ330ii1mzZizBphnilUaJ
fc93o4ZneIpaO5UZ3z3htNRF1QUhwVVtq24bkbMoRAMG+CilczC2pNzirh+rLJ0oQYXZnsK2sa5u
CK9NdpCa3JfufBgz7arUmipsqxrBbZRZ66FyyAJjoI77SmAhXR/IiVyW8ANWKq4NfAg6r14qa/wI
ur/A67mWRNO0N6GrKtmMz6vXwV7INfSUEgHCm47fSykiDV6chE7gSjKe3axe94eLE6n3xd+mU2Ho
jJ0atrq4q/5diBy/tnYCLV4+wVqfQ8rBeWlv8eqM5JyaJbuC6k6CWG7AK5czIjUjsivmhTxxIEY+
SMTdiXL4XyOkqg1gnrzCw0+1eHUTELU5fALz+OJ6lh3Msenprl5IID5Y0mG24N9pXSaMlgIh11LE
YKr2xBeXDRz8J4yTVG84XfIECYTdgUcmZLahSv6glltyMKC6pHIcg/6D0LLKH/l6qBDGMU9NifQm
H+O5CnGRoGKdsumP76j4sWmPIvTG+vNHcp3evh0nwnCGDdwuIh1OTH8gTn4gehSGaW/X1VdHZ0ko
563z9IH7loIGMGGWMmhHG/upb0kESHuEHd1m/heuOsyzUp3DIKn+4+HlvMRXjx8YyAQK3eAZ4itX
rlalMbkZ7QV05jwnJbhaa3X3zMTG1PvrhK5l+u8Psau0ms4hZ0VXjjXVtFEAjTH1IYWRq+Wx0bzA
SaUf/hz3ej/BZPfhFT1zeEZqzOoHjcbbcC7LivT6PzW9gYgxheZj/DtPLAehIvNepiUp7yFVuXaR
FQ9OCu/Jc6QpNznkGNdUU6T+pA3O365hyZN20gDWwGyvR2/wuLgvoGf9GO6vpoQKdqAZJ0BshXzP
hFocLLtBUqS467ROXFvqFB/X6dL4b0BcVQSvidbicLG9gn+H3shIRJJ6LVuu88nvblVBPnAbuW3b
lbesrDxxZa8gJ6mlzaI7fDVqaSu3q0JY9cGxVrrA+TTN8HX9+rL+dHqyv5cGjoHUTS2aGtMOUAVs
IxW/Kz/U/TEwep4I0fwMFWBaVULKZQ9JCEHU7hSNpuokwxgijldplAPEk2C+bVNfpS/ZJ52S4Ayd
PIZ33CeuYfQQyZa4FziVHkh0RRjcRgtWatZXWtJNKg8qUwgCC9/jdc6K05Vlu852Qun1LrAn5WRe
+d7YY9NiSL70S6rB1gExMcEG3c0xVR4iusUvCJVW6P3fCm0uQyVoM8cPKSVw0Wy8eJ4Xh3v7braZ
k1YAjQZDAhnCCPVxwiYQWguLjqoauwYg6T+eGUMcdK+FS3HEkOixXSljRV3xkTbhUGwrCY1VLx66
cP/4XgxR69Zd+RmBsL5Lpiqp7oSbRo21nqwnSF0Oi8aUhq2Gquk5rDo4MMH+cOFs1dpabfc9Gyb1
XMm5HVgIgVhMjclLlOPfP3+0ilw7c1OD8JvgEMna6ASa0hw/I7uhirSy5dyjgh1vMeaQQSR4yewP
PxhI7vEbzFCnbCeCfLiXt2UT3co+5MGMApwRga78bL/TUAD4hgUDLo7ijA63sidnf+3RP1YiYmr8
cap36hPeNAIlBah9qNvBBLx8AoEhWW3yAyFtlu8CxoBvpa2P8ZDkuxO+BIEXk/6SLpV5vGFSoEcn
we4KXZQxQPqyV7cpkMCFDeEziM5NFgqSdBY+BifAK/RyLww7RkIxivLxZq/v/oiafEWLr7e5xcJ7
6wOH2x1UFc91dkgifinPqJm0bQCjr6Hr8/IJaJxDUJuHMIPwli5dmG08ebtL7xXEQU10fVE7bgbC
CB7koG++rs0KOhd+CwdYrFmRVnUM67M6P68ia6nV8mjGFH6XDgHWIzTH5sykHcw9pmxD9H5pNCPZ
+urghlz9xcwqw3sIDri6dspEpVVusllBt+dA+yJrDAkwKm+N9ZZ8k5d6y74GoFvortrTgtbXsYHe
ZRuU19wXw1UpK4vZgP8a3rBDgBBm/YVuPErCXkHlk2eqUEufoeutfeEnck6I7Fmqn2qw4bHxbTaT
0ZrZvH9ezq2xxD/YTyzNCbkvJcHqk5J48fgIDwNMAEf1PgjNx2SIY9SYXMxSZkNI/yZ7LJdcNrUq
vwgzcflY8gpidMrP7OXiPXUvNcSrfOXgnCAxgcHihp8gRTMDDVlReOQPghynzOovYTHQCCnvDr8/
hYChHvoKQb4vAbZPP2Ny97AYNgBVVZqwdodFX86+VpEwvtm1PWc+gzF0oCGNJ/MLnIhdB1YxlnIq
VdNyBwy4u4XTfW0Nvtv2oizhSUE+jXxGN2XYCShyT4w0xvh9MuU+G+fCFlGANL8S71AejWWd0pfA
Z9FWw2xvP525YGJeuaBhbUC/aloKNRB/t/olhfiiJItSqzOm/H7XyRactQfWkrsvRHux61H2hTcy
j1OniZNBZKZGkHGfr53FR6q/0m+CuuqlBYq6BCWL/B1Xa4hDmqsCTVDxviTQ/hginvEbEibApW3c
9Xcwz+pLMU2vBI9riaUJ9dy5yahW8xtBkm8SofmO6YFNBlcSshBAWUkCda+100K6QUGqFX6kfYrZ
j8il2gkAxq6wYjig+AvfnGgI2m/a1cYDLCJ1BKBVy4NLNIllA5TilHjH+Ug3jZJwy6hCajLx/jc7
xCs9enIyisCOtOHFlUWgPbiqHk8QxKLBCmhubVDcWlucGfzAqylBrk7jUC1xQFUvSLtnm9sUTEU4
st60n7rYZMTU1I74npvDapKteMETlWtst/GJ3Rw45S83cK84QqxCtPblcIaSzl8eFF8on+2IZpP1
8bSs5ZppzQd2WMDnW92puHP3dPPecwgU1TMMfeafwwmkmx0hY6W7x6gq5HgcDSvk08VSmmSG5TzP
M09EPj6YFykUcQXEkn75ehHAe98pATuOQP4k7sAbZYSrYt1mYUa1hcGtPEOCFefIU2qN2IYSy3ed
TfIrZoCYbIpZ8p5A3M314d6i7PguB4F6XwDxRQCsxvxxjQrxFWP+flvGytsWmcKNVwzpFfB/6eSF
Z9ruaHaRUsLHJW/NrbG7ifeFTG441lB7p9WlbHjPY7RPhqnbc0ISPpCxRHnmOGUl9F02PhjKDqX8
XzMF0LRvJPp7v/xMp8jnYsgiXJ9lI3bWHBFfrOEDV4WYGKQw1R4tCiMrKkyu6tOZVRdI/OgIsjQH
eEUUTGhLecBrjLhkpD0Zjly1y/9a+WOt+9VYIRkw2lm9oEhPTrrnrTq51fs04gIRCKtT9wj6/s+f
7QYHaO8XQufHnSF/YL1dtY55HwaEO4zwJQ9eXXZD3LOn0p/nuqesqTipZnufuvAse80ICW1rtYjw
5zn4vCI8bImcpx/kCgEUTgTQATkVypJZsukLYTqQrJSbVgA8mevps6cw+WpK6YaythhDqfPZusl7
ljRezl2Wc7OCkrZWj97t0aRWY3GEDdA3sRn5S93yYVNohEJ7KZ9RtMWsfUem6IVkr2YoyAdeGZai
PZNpAN9dSmEgGGr057w43fHtulgJTAw1fn1LqGLF0AGnv0emN+WKM9W5Bid9TgSpuaSUcYbF/Qnl
tYZ2hSJU4X1HUOaoVVpCaggsZfYoqTGMAia335XNxtCSxOBKRUUU3e7wxi0mQKgC2VY35clx1yZF
oOdbQBzgRBZMdLEmuVmTS4Vr9Ww5MnEwSZwTY/Xc9qUM/Momqg21HxTpT+7apz6yNxI/SuOtw9v1
7w1vrMg2TuOlRO891QjHylvLh8LipDNtcVJlW3KUQDChJMpB2hUWEyU5ExF2Nv7BYMUu4b+mQo31
yvP2qr1cIr044RFxkMavVQt5octXtN0a/+R9Q3K0kxNQ8q4wP3v+jmebTj/92QEQrcIARg20THO9
gjboplDjHCxYyeneD5rBy+khK5eA8qGVcTRG51sDgcNsAM5mbzBsr42PoXh1IWTE6PVb2V4pfXKj
Na7eEqa0EanIKfv+NiYyu8DetwLpqhf+7uboDbyvoy55QEEh4I13OAkTiZskJwNVG2uEoftuC2J+
COrF154c5WkSMb6eBD39XJMUUIcFb3Lx9rtoSpniPH+LnVLKdDei83XvBSoxvlVL9/qZFg9foN2L
YUgbJIuMZtnMl1j4N09heQ+AqiPexNCOqeyAg4O8SohmjstXoOm0rmY3UPSrWb2crXLWhIf226bq
7pfkViiNAgUSiQH27xPBeYbA05xM4LDFuIwHGx1T753p1y1/44cqurieYoNwsEhiXiycN3pHjeOP
lLC3QHhQR97E18thVPkkl9p2O1BMj3MZLIm2t0uAI1QujhuCm+M+uHrV/JTdzCJaY87CIgEnB4p4
tijcdD6/eu9mAfpuBoiJpI2CEsSnlueRUb6oPB7qOMII2yl7hU3n7EzkGOvTrMAPjVfoSX3ZzABf
t2xwAP9MpIi5Zzx3tvtZkegSdSw6OqTwEgESmV7n7l9sxJwDGIYTm+qijvDcgT3kbG5tvr/if1n7
l5+r92ceoJIB+4NBupsZMtlKOSELr2mB5sCtw6E/dh4mAhQ6f5BUpVJxyqLk0oHzpOCKdGHoCmDt
0fx+fpBGr6yonhPGXZvCjinfjlr37VqDO3thoeM/3YvER942OQAGqnmydepcGaGI6Lj2XzyZNkxw
h54ztnWgfst4o+sp6Iyt+hS0VbeK5/WC0RHtLoLug9EwtX4J0JykJjkYCzFFfYtt2tAKtJo2iL8V
NnAbJ0mU0wP14gazjFSzZGdBLABSsF762TCyZnyt5HN7IZXG6O0uK4pcF/LtsaDiQP8YeeovfHVF
1Lhe0xjXZiZTxzGFLp1TC0FpeVcsFin2EUGOo63+lBOZqvG5MZtSlGqUrntgiJwE05NYaSQRNEoz
YJSoXu7S7yde36VDcZWcm0A5E3SHDN0nnyLqAdXoKMmdynZtNbzDu3JKvAF1Hh/S06h1bdAk2lDG
Kk6+zOWACjFlx1m9oeLDINE7xGTFjkLzCw24PxdlhC+dYB4510DEdMLKQhbW0qJyOc9jV+CK1z4p
UYYeWk4OPr2RPfVTE4FvI7FMp6A/Qf5Pfr1N5fCYNmSnWEs3Ry7j2e8H2IUKPqZooj4BM04eJhKk
E90e3Hr3cwJog+GsYVcnV5SZmVONklWME1PsTwP1Uonb4aHkyTceuluXrhM4hsOAHQUuIyaqbjsV
jxLp6/oTBMeWTQtQxhjQ5PqBHkYwh0j4BXl18ZTIVJ3+Wm+IrXtQb8A3Uk9zMEK9bSQ+yB8YY07O
yiTJI7vo/CQsZAGNnJM1GVPGwBj1K4bNG+Tn5jSOdKdlnDw9Z9fT2uggQVnOnpETNdjLWPqvIDKZ
WD4Bu2FukFMa2YV7bX5JWZ5+7cE7AKdOHfuHPEvypiGqChsWRIRpSIcm5wJwemzgM/jtry6GpPfF
Uj/vpSDiGt+OlcSCH5FlDtWUXoYLeAlGYswvu5kMzTXPTpL0Lwd6KFxwgKJkw1JuT0pI0kfaQwkt
sXJRtSVNnMVp/UlEKQ83aUu28UAxi8+dCHcN7jcIAAaCR9WmkAHmMp2L2k9AWnF5hNij7xrfbDxs
n1r2M6UsOk8vCKGduI0J6jhQEZkOYwku41iNkQUBMOOuGIgKRSgjXEL6q4xUjXncq1+WXeCRqpep
F/WUpft7jO/gaTb4mGztAOCGDjtPwp/oBzHCrgTEGeeQWXYZ5hqhGyBk+gsOXLGmz2io39GU3SxK
+tUVgoQctj3Pf7i1Arwz/WxqPvmnHrw8YFO2sRAk/bPgWXj5QVp436DpkPB3+bb91+v+FazMsclR
7Q40ccv3tG+viOCyiKtJkQ2Dj3ySOSPLITEYLZU4orTRfgkrOvq8aDFwdapdMp2quo6TDcR2c2X3
69b5VVEyYR72YvR8YMxR+4uf4J0A4Gf+x/PuCJuzAguznU/yZbetGbJdW4tgMgPzRtrr0qSYgKIU
iQfNooLIXIyvoI2vjLbJw+M3+i5JXFHO9Qz6tLi2EEr1lLn2Ea1OBo6AMzvXljKhhNNB9UWGdbys
xlJLqfPWWaHmnd94vjLmgDexFPy+KwMSgTsza/ATmk/fDDKP5JP+iOUUXRcsvow6LItiySilIDGe
/+WayKKNtyioLOwvi9NH8NG+9dZqBsdWngIVvvQv0s8aVtdxCurJjdmFMlzSULUstUoQvQa2bM2w
MURpbBCW9fK34hsHD2EYWf5uI3cyMfpdpfo73XH82kozpv/JhcOR4omdim3cdw2DPcDq9Vr+7e/F
/2+/2MPwEIpmaJk9a5XbooXAgeFSHntM65l/2LPMmeOTfIVPhKYm7ArVx1u7Ig9EYnXj2bRFkkYi
MqCmV2q7+ulPrHeIq04b6hjiqpaA9k1ASaL/jgWo7XhG+axEq83ktCuuV1HziaFbmGhh3iHg7GsB
d3GalBazBUOxsf6WubUDxcbpyjTLrOuHcsDyjGbz9vj1D9OImsbPsGmHSS/cQuvm8VTEu0ET9lps
p5LOm3riTLSZr8thri/nvtPxfdZfo0Lyc1q9/kSMWDmNMte9QPwTikp+cBiHZNCOzdW0/YpJTTaq
MLeTfBV1Ui7gw/n/79WDSH94PufhB8ppUp6Pr3SW0NETJm2OCbEl1V11nvOVGxzPhAIGgr7vacVa
FVPGm6uN0fBWY02CC5Q7+kohebGqotcapkuzdUgUQ+79GP5LAC83hlcxmD2/R540gDO9AkvspNL1
HPqAS1IjLQBjJeO/v3XgxByJI2AIm1Cn5stfPqE2JGjCZ6LPhfRZILSvwSKD5touScf/N8MPg3qe
bAWvIordrv6ibm0BGc5gNjGqNmHdRCrIim5iV5xz7WACXIIdpfLhPE5ljcpMM4AetQujw7FGilwI
56PX8JdRCh3N5tXJ7/uDf4UcEXAUV9v8sgzyVsiP1mrZCbVrwT503cmmyjMvhIy48gL/BNHIt8VQ
TIJwDRsBC9f9PBGLZ9txphMS+2E8ww0za3lwegVq4z6huAaQ8xDv+c51tUTzv5P1XQVg2Wmjiy8j
E/3ZaT6KJ0hBFmGMz81vSXPEDSOy2/cNO7dyJGD7fdt4BDWrkVKfL9gpEa62elnJHjwnVvlU3po9
f8d4ezKFb1agTh9r9SFmu26BlAqHFIauefFJyoMbeiLOUnRnAC29DXDlxNFYNtDhyN3+bSzyMP9T
o7520mQYuOHvwd3sFtXAaMTunhu960bHrXZqqKWdOqobG51LDCS1IOpbIVyv4+kDz5pDI+W9WF0X
bHqG2OlIg9Dj5ZrKENeya8PZedO3MVqXSu203dg/FIVjGzas7yScfPeMpDV75ka2txMTMboXE8aZ
usQcBbuVhIrtNpKe0xT7BNBn6IqNfP3CMNGKlgQJambPlv3jtBozfzlqwaVyEeSBu3/PnOaIp1ue
qrhumt5O5DgNxjX5Lv7Cp6eYmbwiH+5+mAcCYbkxtouzlYcGGv7KILJQvGQx9jUwVKO/QHw3yU9Q
SHfDInKaO8mJ+sBYWZ4p+XbD54s3rklRnUJHjrn4x1QXGmwOxbCZeuBLSYRMR0XYAdL0Ezj48MDw
HlL9R/651UkzCLRbk630BcUh+hqOpEvfMcxtZ581+s8ca2D0eiN5uX1ZpJ+KX8S8OgJuqHYaxpUz
I/97t4oS72hCSm3omx5Kzw4SE9DgZTnMwliggcTkIGQtHqJ9M+av6qIck0PTzAeGhrOaHVBm5vfv
cEFgTtYwicIWIyYu4Pday3YPW3qk3wRLFCUzrR9Xqib9rfFqdG0A965Q6Q2HTlJ2vis8EseO+Tbs
tFy2pMOHnAXxTvzoN361bGycr3K03CRklJsdWclmQmJIsGynD1hkei7g9yCUSHmEK3t/wljrtW9/
ko16Maxk9w4XFDYV+jhFCNSPWjTivBIYvw+AiYS8x1OFW4ZNcrAqKKs5790TZP846pHb6gGzKi0E
9NITQVMfRPyYVDZO/pt/492lt12Py0WaYRMR/6nKa3yhEYo8hhcix03kiK1FBbD+sjK3BBhI2WPG
OzNXBCQRlNzGIpEA5PKuJOhrmhZq72iUhHIg9y4M53i42bZwAQ0ORyFwkOKCc/tiyDUtqmp4t8ON
li2zzEipO9u32qgnP1Br1sKQxv76ZpeWFKJ6e2qFxZdmu19O8VBxPntQLuKYAwoAqLgrhkvQhlNX
H+EnE/becfWxMhOyAw9Apf8HpW77J5JKZcKNB/FaYjfLY9pNVhXzS3DVP6XbEDgmn5AvDGJK7SlQ
UHQoH11j9s0hwSHRsdzRLEw13Zj8K4CUkixz7pm0Caj9CjsnuB4M2CFZl8lqCP5b6pwM8lIY3fhQ
1G20k/g/Bl9VKwJnQ0lXMqgfbuq5+lgiK9RPJu0WIMsSPF6uFV4ytIB93SHbuu31XvYNu1St6bvi
t0hfgu1v1TeJPP3wIh1XeaRrPeKQxYQUubC7gtLmHr88EQcJerXYiywugkX7U5KuqJWN2uOBi+H1
1ywbcgc57/gRd1F/dQeO/qf2FE2NjAyI0ubxvt66us87PtV6MW1RtwNpmnGn9AkAifLiq3zBcR2W
sXVsr+5fpq2iOOpZ41LxDzdwtSLZT7Wo1roRFuzcS9FCPD6IkIj/tQ0OR2Jmcdcmk2+bnlqxSJ8+
zymwm5WYft+4KCKhuqkw+bFqDPX9/lVJ7glKbJBWsMpS4gn4q/A3VBKnrka1jtPlRamXwK0U4C4U
69pFhjhkWjMeJ6nSfAO9Jh6fzUykRe6CQ/V+dSU28S5YLANvnB0J1k1lbgiPomWGhovX1cBm48PB
MQG7MrRknp2KuS26Cbar/U8EceGXEZKSDlYWmQxe1LXsd7jH9VeoEzGZGaJIY8JeshgFi8C0jlTc
tXp+78fM86cHYt3SjU9WLBI4tn7Zf3FYBG2SuI5fnJNahC4ZJU9RX1V7dANRKDxiS1JVlP0Fa5Oh
lfiiAuthQ9n9CQWqOFTXWLTkiKr/a3rV/Qyn3zMLd6vUZ+3193sXQnplETxWP+1SR+l7+yzMbLwl
Xv4T572xDEk5jmgTfVziwMO+F8yFH1n8dBdyPVtqt0luRBNFFjdhwOvZ9CbEHCFPgpDXTiyjNx8l
vhnLXSiVhhOgOQtHm+grnl8Bz8TO6kfGW/LHJUXL/vM3RjXR2Y1kuj8fBmZC+t4iKnBSscbRDVRK
O+1Awtdq3Z8gFqAWxvC+RPP4Fx6ocw8+5pWssdVZnL0wZQDBQglckuYFAo8ZoC5BkrKZowOgCfGD
etHpvjzhQiUgpCeNkhZfsxFMSl0iGITZYhHI31vPMyoDCLN3VF87vbIPbSp5uh8xHTKj4ck2bxci
yQuc/f4nIqTl63ptcC2PQO6TZ3pVr64pk0dRfXUcHT9eQuTRa95Mv9rPjN123vW1CWFdxljFk1DP
AWBGYhdPAKygPpALBFCjCm9qsCGZalfLeFD9epqI7pyEzKoQYaVnSd9P1S/FUTk67dh9G4G7UrHZ
v3SUJM4gVgLbcBGN3fU90ly/ElRGyHeARmObv2+vXPJHs9wUdzP4B9F2QptqxFuKtjbZ6bBANxJL
BYDX9ENqMg/Jn8muBO2k35+b/aom+FrY2z/Pw9bMl3Pt53+vXTkeU0jTuC+ZexhMhJgFmRrxM7S3
tJp1xuQ8XqaKL96uYIDWmob9flDYua3UF6ELTnbGm6VOYsgU5E80ii1rJYRErhfkkMuhwvtLpIoy
YcbZfOhtUpQj7tgJWlVu0aKA+dAS1PXckJjSjykxpJyIo/mR9cLbJLtIW9ZmsSzXNWLo9fnN2bYs
oQKVpuvnEmjP9nPi8KWc/P0Tur5zgiLR62zB6GywTkVu5Y5ymSeW0YX8sm8AXI33+ya3nNFsw9hF
UJCxG5YJs4vKevuePlcgyxAiYhPa+tRpJWIl+/b7/eqR/wB0kyig+RubjN3vgSyTiva1c5rAgM+w
b5b90muGxYFYB4pxqRMZ7qeGjvQaEFKt5eo+XIxmnut0iAXSzwJxOtDaIyNN2ON2/qXmLHcssOJi
5pgxEf0zPuDPBBXC+VMKtkUwvS9yh4buPo74ZdHUHhIJsbkKnYV0fmdYK/09UbSHVlT3EQhwlgES
Uk2jODXoX6NHWC9voTEatoC88fnwUROnw0ijbjjDj2Vt9nsCH7NBTseRI1L2YD+f0cCY6Nt1aArF
ACjQPVnwz4tIMjWMYTvNo2nNUrZBXAgmaVcdjbOT9RC++2EwhXIz1JcGPkXKzOTvO3lGAAyKEDKh
q5GH35DkFf3qXpoIJqLUMA+SzCmvsDQ8nldwQv2TY9v+XDXcPKwlh+M8Z1mT//0+DjNDJVf7ZOX8
ucTjHY2rcZTXBW1u49wR/rBI/TtOArzvXAGjAEjrQ96hCles/fhKlKUJ3l4jAbCn3s+DK5/6AJ+E
anjVHAp3zRPYt1Sl1nItoAN06l5du7NwMhLid9/GZghBwI/idH7//UttaTYzEV38Ocgyicjbpi+M
mnu7oqdcEWF8Dtd8LsEMpru4l1g7bQp/hal3TBWjFjNlhfw8AeNUXN7Ref+Yy2iNozZUs2fuHNGn
AMhzssge/S8HAqm6or51eyFN1akVO2Zl7c/hB+9gwN5aJRPRJdAOXC6+60hRY37LL7JjlAwJDtZ3
FXCVp50VEgJMXomNsF5yLbwoAmyXL32sehsFf4umFbaqsVncb3hFQ9m3zJnjLr+Q8Dz0KvON3qvb
hce9nQnXJaNd8xpENIgCsa+LkxjLkXeb4v8PZCKBMGIAB6955oKkaX26X3BzdgDtErZHdXqr1FdQ
k3F9iIdKlO1gG6BLJgryKJtRAsL9hKByv/Icuzf6u/G+5u8TBJdzcimsefycPnQG+4gd223ixajH
TIJZ3p7SGSoayBpSzLwngYR+4AfIKFumXFl+qxkIMyhjxKwpSLZG0Zzjj6wcRLXyhf7vxfflC6EE
cBA+IipOhU1sfwDwZg6GGah1QGDFCz9YaMlSp/IhBjAzRhtuE7ZcrKk2uXLC0EnI2v1vLVV15iQX
TQBGbYdw9cVxa3uOHfYcd33ID6w04YCz264q2cMpcEJUUpzyX83bG7z9NAxFwXxv98ue7BcsDlUM
7QeEo99DRZFhuv2aA2cUu5aoHQekiiW8SKVxQYYkeLf8+4BvFEJP40itwfh0Y0X7xtwP97g0ms2U
f9vshkNdAZHARMtoTvbAzg1+Y6S00WhDYRap573A3vFJ7ku9bopm0HUKzfSNGsdF6r5nMzNa+sbt
vQ+BFL/pZaaxfL/G3+6qH/+k6aDCjToV59qrrIYPKcEMC0sd+o9Daxp6c+L4BB94Wmz5M3dHleJr
go3AAdXqfrILtI13tG0dTOmXGa7DiJR/xlbPv3iafbbCmYgFqOYk63DUxcWAd5YC7mBU/24PBHo4
GKJQqREHMVaBoPkhVAgtwzrLMFLNAVeWWLELwHrhvlZQsoEBFBFcSfI5e6EhQSANaKTYW+0TfNME
UqIcD0Y57u3E6UhEc6J9J8JaG/1b7WohY4h54ohaUITlulfkDyXDcfREjikEIMKZh1dwrYkqJO9W
7Xl95F/Zx5yugdy+CjWe/VPmei9Tk0POQOIXcA6YnqDOb6SFtaPI9nxQz+0weec78bLFwUJSX+Zo
9qUgCJ0vjBtyRGrxL5R1UbiiXj6j0Cw89Vlh9l72rPoZ4lKdbbO7ajx5AGi6p+yXvPFXmqEOEatg
t7gTceO/K2HuBDSI4IusY4tgd2f1z1ZGnCqY5diw337U8RzlgnWmwaE5aFnBSxxlwdgU3TiBRxiw
aHDB9KQC1HHC60JUWJIU4balx2enW6tBnOu72UunHb8jtLWVfc1CPYG99zgLVucvcK8UwColn02n
vCtDYsCTmI+R2tO6tcytGx2gmnVQQNK8J7zqvWlJy9ha1Ecq5lR4dWJ2xllLzjarWCxvMZAFoiWN
uE9OAa/5cdmKksJjitaibcTXY1ebsk3WnqiwqLEQJJRJZMxXWQmWkw4CiAwXAkulEju8kgDTsUEE
kmFQ4ShnYpVPzmxisMboNJh7XXcGQElu5Zi8EqEIbhEl4Pdd6E6iry1QWhlCUZVTG2VR4FxKlP6Y
evBupQem0WCsD3QZgwpQwIZy7kgpcB6sn5pdTclAoJZQUjW4dAj2uzUe9bSyOwLGdvu3exvwdhy6
yLHOkiBHOuABgc8UbuSYgLyZxINj7tsrgdx2CovaajMWeYmv3j2/SciRmJqQcL/P7jxBmjDvz/Gj
9qyXDjYHxMNFDPHqB6I7e+tw1832bC8flU3FNKhyWxTrndlvdF9uS5kVciqTSLKxS/AbQ459NSJt
FSLHWi9+1+ygUm9m2pmOHUHmIp4i+92KGU55PyiAgXi9uRzzFxZ5xuHdQ4f+ktJms4aP92/p6/KP
M4pfeE5GZL0sOy7HuQGndtpt3YCfXVqgoZbzk84t4ZjNCkRIdvqpxG51i9fi8bK557WNpjMSgr4n
DtI46CO3YzCZbWgt7YizJfnhnfRQja0quol+TZjCYm+USCAIH4kLT9e9lZCHaRNMMkuyy0MbAuM4
84QEqvFPkOX4pA0rwsihuXke3wOy4VNnfhA/hhko/cVVqG6MD8QIEzQ6ariG+6QJPdgZVBveUwRs
21StLD5FWOHd+9OTGTQRvOP3dnkr8Hu2G0Z3zmv02yLY9JRbRvHsqYvvRNnu2pKL1xEITxSaGKIP
2NTkZom261L/gyPDlERtCkkcnhwtpjCY6M5uqn3CLQtGvW8kRt36FK1bDi6k+tlCbi68XQUQlgR/
Bgjj9IC+330y/MLYYREnG2VxwOeATm2Go5MTnY1YH6YOnQPrrjY51zUPrfD3hio4oWFhq7sEq//r
/efJR25oCPN/1u3na/4oz5JFArWs3tpLCp306lYH+GUXmFC5J2trGJPkJCkGM6htPfoFNRC2Gq50
hBQKbEbaaaaAe2twAXzYvXBHSJY0UVJgyssALFtGHKEZzUp6RrqW0ecfyjid4QS8C1Z9tyzsHSxQ
795RKAxbWdAYHSJuwpryv6DibnjHfOA3ND9CUFw4Mt3qrWMvwufTon8tHrzkVLnnVO/Q1NhI7MzG
L8lDl5NKBRGVkTcjjoCZ3s6fcdqjNeyZMwI7XUuIaLiFO6lgrAxXGZ3LDwPdaFeg2zTvh2sEP4j+
tkxuCqOhr834nhhlQbGa5zLnloCtl2CsUROSKtCXoX9mBoHZ5swj/dNO+nD+b65ATQPaZbQIzzp4
ypgfckJfBjWY6JqTWJ98OqBSThy7o7o2P/fToUFXMeSZbKNo8ClIzpTXzOrxC0nfFQpJk9eh8giQ
do+FX6UPBlCQNbDVLyGFc/gtrmRM9lafiDnzsUJQu081Z6HZTGu+QTzQzfrrRGINxMH5cSS5V1O5
ZNP77piHmOBSpPgtBVBwcJqcZB2ukN/IOrZLJ6AYBi+7A2IJUVVXGGX5Ftgkyx9iYAG7RfW6OBr0
W9gVWUTbbGmx+oYmlYTOy1KEpwGyKzcbnw+HvWqj7e0/whiuoGy9qIxFZJJ61ASFxOQ97FuNE+dO
K/B0bD7e/Gna+wSDofbVjiSjKMNO73FS5XJrcbFRHvcrolfRnBRW8chUyNZe7rCPRllOfWG6fGiL
D0wiigoo/CkIN1taCDA84EVAq1dvNXwoogPbUoSJFzJwMmElAeloV+jWmzZ8FMfLn0agK+qksL0i
yEGb/D3fp9+EUUDHT82J7an8FZiJBD7OyciQulXMCCN9nHi7DHGYwJPP5wNHfy1SLGOAsdr+HLyb
7BTiF9lwrrFAaczUA0UXydHbPAvaPD5Mow391peek8C0Ly2chsKmX2j/aCauLa0HvNk/sgNqu2V8
sQK5w5Thl9UCYkP9wsYbSpYu1ZpANxy+DwmaRl0U6gJJDPT+qLkkesAYkHXbRHQxuM4olIlEOM6S
sMOdLaTbMecs1KIPnq8v/B9hbPGkeMSgNrUJ2nFlpe7Jo1esKqkLjpfPmN4yuNoo0KLa1PJ+LCOk
AWUpUocoPsH6ovytXeKMrtXbOsa7244k5lvqeylwcN6UuzQ+BUW9/RdN1lUcH0aXdDC3I4t/pjHc
81pfuVLJpl0puCJwd8ZqOX9RJgrXmubEJFkAs42qQjznakTudsBdxiAwz80MTREiXCFQDy+VCznW
JsVqPbgdayFRCSRFk9OWKnQtkGeUF2R5VBxt9B57+e6jJiQBzcqZoF9e49ZsLXWfrTa5zU/VxGcY
fSyTr8vZq7RFWeKkV76mKSdzGBOWY+K6ZrOSc60Hc+yyXXK1+urEvmJDD6G/qVHHMJYvEAYtvoTz
F/RJCgf+L88pRwli0US/KIyPOPd7FiwUIHW1ttIBotop1UaDIrq0SGahWuDDGb88Mxb4FFiCUON+
ApbcTTU+h2qrQ7fgi5CwcfOrCXEFf15v0ilZM6PknOpWc54s0XTxyI9pY7Go9T0HC1F+Oxd8tOei
1Mz2BOcE2QRj9Pr99bSB3U/E5tQSktwdoFzCO0/3tpSCi4W96EV9fpltSJjDkMyoLY5KOEvgDdMq
eyzs4rI1R6tZkUewSYq1uFK2P27zF7O7pOEmD6B4gMMDvd2ktAfMF52fiaWQlOBWlHtuLxhXL9S2
KiSupc3VKb2Ea7+AoUDqGgoEKpigBuZuADJbWd6dCqKR5OlR/dKD/HJTzEkrSUuz4+6KVBgnfm7J
k7vLbRTZn9tGaDuvMKwQ0Wo9ryLIg7tu+MroMbe5gK34pzoIEdqQiJOfoDH9okSRlQfuXX8tYMXC
Bq6cUyLNGqBguuKdjFvHfjAWSW+f97Z+EpDfYi42laSz2twKRQB/9iz02dXxSvnSz3d4M4uCtclr
W6PShK6TT1E8Yk2/P//35yM7lbgHdzfiUW9KmCL7ciVdtsWfcRxoz7+cawAnFXCxemZryFPIaSHG
QnDFhG7jYORVk3Ako/jx1EKZ7EeriluxQVpm8f1l4h63l8iiEKE92Zji/aCwp7u0/XYi37gP/ApX
cYCA0heONfonz5mN6Tv1ChJJ4CbP6h4kDOEjm7tlPWOwJeeCYlAyPAsgNXif4mqxkv6UG9IuZw9t
iRCIvfkWgeRCQgRCJias7Wf3hxTOOjlUidDz53BObM2zo18BJQw4CR8z8emrlOkP4AdMbHJu7shE
mmXu1toiebJnTMxX/LhkD3d4+0wnUOW863FIBqmT2Bg/bWSwAJPcPkKQ0lkJY01rmvzmscufaM4x
baTz7mTk4yCaatokN8NyLngvFtokxIwCO+uwz2n/RdDlwT3y7XPoGr9Sh/NedVjswEjO7kh4HAdN
ISCGO4pnEr7jClZCWBxFBqxglNglP9PthBbIVqOwQ2WeSUKeNbX0C0WjW97whkOCWjXsKGiByGLh
g64wqvxYldhSLyM5PRkg7lbgnu9W88i5H2yho7gpLWQlYRULnuprSrcfmfE+Y6m3YeOZzXnGSOps
tioSyLjw/xZROLYEnsbjVEQuWm9dec4eZBep65AI4so3jujhI7QXcFCui1JJmU8HWAJRzM6lmBnm
9K+u+NhkRMCkId0SJZUilmdb3Fs+1rq/otz2r6obnVNe+5yApAJmXfDlRDeFNRAUzAE+DOGvVYCh
GyAyQrJsPmd9ZZVt9qW23PHe/dlkRvwUwNWlPkoHIkPALpvv56U162gTQ0Jlmp5+KFSZ3IncWBqx
hq+31oX7BDOUi1gm/sdQc9+MYMODl0asXfxexUR1q7V9MJwyyixuCSio2khfVc6FGbeeyInSdbRQ
Pztyr+Pdp7Es6rOy2iyBgSJErYDn75UqH7BiwK7jqNa1T2OEC9CXH5N/AdNrFIGmK/ukaGDa+ARh
9edCr0HV9kDj53rsF/XNCWUGkBYqf7dApRynfJt+78A9vG7wtUGnJPx/3b+QK6GF8CbtaeG1gjux
7vRiNPNjODA69kYCY6Io9JIW/Ee1RD0t/q5qMP8++LELgLCZHX9czaDY15j656H/UbKY26V7Ttm4
+0JxtgGK926XDU2IoH9USAeedlp0QhC8OIrHIyAEB7fG7d9PmGCYRnMe3aQDnAOxecqAfju41421
HHjCycwRWL4sbN0jl6bpNIxowfO1uZ0Jum76oB73UEOamGc6XzIc11n5ForRK7rmezxl5Wy7EMvA
KSsXt2qHWh1LBzjWzGYL1Is91Eh3wXlVA9euAW/fG/n0Jk5p5iFsZC/6yxSBeKmwAJNe3tm6TT8I
54NyUebHEjCepnLbrwWZ0kxYK2rv0ApxS28B3ihzzFxEmqnGh37DE6wT9ApzBnl36+I1CJttPf/k
KR0yLE6oKdmMYqqjHYUQW0BPEMrgqBZEYbfEcuj00EikWNBNv2xoymCUxjn76+KWstR4ZK29tupe
ejTLBYVS81rjNGhR7QPTPJOb527zbb0QbFyFuKgj53pVGY5v8fxekLd+G+SE7JCGwfWTvJrtjgd5
7nG7VF+aCnMtIUcN9DNh82WRCwzl0V2V+VOdjcqqtkgfiNQvqwnMDpoVjxbpnBxJ47wsH4vqecQJ
wODN9s8P28bpLOZVTJ4Bdm+Rn5n/xUlS5BVDeb2c06yXEONcNYjVsGa8YkuczH23nnmWzoYQ5qoD
4Dvi1cKLy0qxepYJ8TctXWf1A6mfkqB0BZAdRDA/Qv4XKAZvWS5WteyuZVWsT55ocA+QtMJ0Se+e
7iqfkxMQT9+fjXacIWe26F0ylkX9RTxxQ2f00O3SGD5IcYzbBnj/PlxPYTw5RKFsj22hNjDn7qgW
CFo7gyg02K7Zo4Nxt/zNNeF7cpM09QeYg3LnoUQo8ffVKf3GvCWLtLrcAtUnF0EZv1v3C2sKXl9q
CUj+lp6gsdZ7Eus9bYGjnEnDxZvEKeCZpyi1q0wlLPcYmMIEUvkxnQkPXNok/Yfk0CVqBgGmvC0O
wF+OS8qrnM2UBOc3BaY+nQ/6GIsC6Ghvk+c7c4b6oJM+Gi894yLauL0oHtJVbhnIK6vIeob1kZII
AE+rEz0+dKAotvmlnCd62gU8BlmeBOXCncI5np4STi3Qbl7Ppiamv9OITA+YdfK0B+65Ccv57ZES
goaZZ8s7HDT48RJTv4sutrnJp/wZ34LBm2gHDQWIkNZsZohfWC0bJfmbagBZtHVC6YXXnvQ3bP3y
MosM2u055cAmR/mb16dGrsF/OEfm+jH8UnyPwfXuMQzQjIsO6XrUi0Sas+170zT3FyQQHMf0DmNc
2KCTh85B9wi24B23uAoEjwMrVXUwQeEAvDvF3mLyB4ymxpwHF3C+kyq1zbnvTEAGLFGforDXbyd1
lw/a3WkZSqcqy9sN1skxk51SM0T41NecuVghFx3bC0f7+uHcez3qVIepmW0bjTHdFppaHpb0/I9l
+bM6GAmTJpe1j65V/+MwJva1sn8dAid+glgi3bAWsG7+xJGtjGkyCj7OlBfDLPJGPtWE32rF+nID
sMJnraOcMCuQ8xw23W69cC0+yLBLn42zUBh2cG6SC/JOEUJ3LW9ljcc17E+3QkvpjJ75MXhPflWK
V8UwQ/Z+nquXjU+r698sOLCSSJfEMYOww67FJ8hefepgN5t57aTm/cYw4dWTLTcqYiwSgmMtDYl4
z6UyuQETwUoA3Ow0BOpCa73U4uXc1wkfcZnFbC6YyHYqH7CjgPaHMj9AMV0vOqT3h/TJPKSVbGh6
QWFlh+dCTIqF98Zzwd6OJOoVoMqLMIkAThsjmIoCBoGBE2uTrdTY4jhAsnCIExDGDv8KcSzaz5hQ
n05WUT4CBD0zOEqLJgXYMM/RNmZwb5ncBhtAg/TR99POZJUi9LTCtbSt/+d30RiONHVuJrwU6KWN
jXkZbIXHB1NSdMKX8ta54pdfykAb7w4bkdn+LslJ7s99/B+n1Upu7mzvj7lNnImJX8eyWJVnb41A
bmyEN3X5v+ZIqD86owFzZ2UdlUaG6JKH5qO34vKIIryJi2MZbQsLhfGwaLQdc052hgbPChmtAJRd
Zh5m7YxipMF/JAf2+yHMnN/HfwOcLbefkjWWofaKusYvC3JImDaMIaLYk+HfAwj2hZE1ck7jB6uK
uw5DRlDc7ymlt/9AENMlDFJFsXpFCmkHaSN2+XAPn9EHKpAGgIXGjHTdvQBQw9nCXO7MmNJNJh9J
X93VFcM4I/0dfZqo/4EvV1VwzSzrMu3bNNG6IB7Cwlad8hYdfTF9MVQjUeRJ4iz8Xw1eTgLydP9t
L5PlePeaEDT0JbylsGrOaCspvjQ46GVcISeom1htHrG6/0iKddi/6+8obEwO/i6DG9jyRFdqQP3o
yq+D9dDWzi/b7GECfgtImjvV2BZSyru+IU3+GRU3lm+MPeRrEE2RUSopKEeomUD4PcjgzHBVEuiz
0kDMZgFCIgP4xAQbahE0HfFYvED67hHGqtXbUWR/CEkS1L+V2mslJvRGAHJ5UnwaR6oiVPBZlHC1
2fknV6C3uKcjNvCPLS/ppJPeMQFMEBvj7THiknHJrxwcvpxja1iEFFKYLq1ghKeMcyGbQar/Docc
wKyQoUjeN1FCLRoJ4+RMhNckdKMQEGzWQ74Mlwq3UItx9XQ4EMSVNWmaWieT7USChi973gZ9Idzm
xy/9aMM3d0gHbaVMaDeWru8QVmMgAxWrHE9sDcZhvvunNxoYAS++BbrPxwNPE8TpFv8Fx8cU/PZq
oNrJ9UOrmi7INT8S5vfRDTfZKbwRfKID6Zy7vkO5zalus5bwdzdguX6eYz1D2EPJGLGDxOUBFQ/p
R42WRrzAN6+bylEULfK6uJ9/GOMVxcDKLoLweGhYOa1ASP5p4SBUxlN3o9GqPSxyJ83CpSEGfw+I
JoprideANJgjHFSIy8DwgoUMnMty3AaIsBLlpY/HQgbUR3ZzwtlsVKPPs3iuWmMq2UKVXCK+aAuM
M2VV/2VzaWM3icj4kUz1wU3gfOiS2IeQEfVFKvlVXTd6l+XZdvUhr3VwuihwZ7cpBZrb0LOWGC9y
D/5KUmMbLgZq8WITidfXBrdxYTC1rij2Ln15y0HDp5GewjgiXXint3NLLcwJOqDs9A5GtprN/hnS
jC2DiBnAS7s47ZSakoVVEU7iXsqN3Tq9VAZExpq8kLSMp6NjGO9dHNwE+KJaIqjgQsxkPsxp1GVC
RMspaqdB6EzzHOxl0/IKJT7jjFidRsRjVao6pQbEAh0QNntDLojNYofCQbCs/wiTHW4AX+4rUGBS
g72B75bSEPJXFgaEpWzkH6S3QGKn86hl9o02sX0TRulTrh3ASXbc7gX4RTs7k5I7SuGJrodQZzy9
+7+sD/Jy5Lcd/EFNnoIpVMFFHHNOcOf9kHEtM89dp2akUKoIDOSd9M680YFLTHZS5ZyRnUjqG7ap
s3+VaWp94F3yz/Y6NhgWizuw8ZtdmzwT0ZeHqvB2wt//xc50OSkm0w/iRpZHmPDeykpOaPI1ixrx
86fWihemlI9xaa0NJpy0gAX4LiB0mXquQO61ZVz02eeo2AwLnffL4aL7AYettCzqDQZdj1L/f+YG
Mk1guCpSEpdgcUsmmpXJ8DNckD6GEJuE914JbtpU72Vx65bN/X7ya02cKmj9Eo4IXbkjl4Mciy4t
wO54bifMTuPk0V4dKhaZylTU6ilzLnf1L0qF7PmP+IZZN1NgEHDJzU5hMVF4TrHx3cJx4r308OT2
+h1AfwlT7tooAtfI2d9Qh/Wti/Mpn3sw9KLGE7wvCMPVwnZ9elFHkHRMc0LsIune69Epsd8CLA+Z
um6M+j9cWXNpNWYzssa2FEESKTzXScSxIS3Maxep0tvu0i6U7oj0Mtj6DvnswWJ6lgzIAm6xzIS5
WlkfAvQnjZxwNwFXSJJfjeqKM5PpqbNZ5VPlBqQR5B/Ru7FHGw6ZAOSR6jJgfPDB+7M0zUQxlgzH
S2q5PBNHqrBaeuSi33Uu3EKIFVMPbLZ52GjyveWulWR/S0H5LNOvBmY1gNlWqtoOnfHG7kSb5OGO
/LmT2Ex5aWAHHUvqV96ogYwr4WbLQ3MpcAKisJOvA+UYAOblX0PGJMBffjJgaXr0SSH5jEfo/egf
JaEtIHPb/aEQf6gMCa5i1y9X6QtAHDjoF+qvIg5DHcNjMmDdUH2h06OXbpWXvBHdxA1fltqE3nQW
o898OsA16+cbvmfvjfC1qxvj+O30J7QGK5Iyow9Yr+jrX61DQegjtN3HGVq8e0Kz05w2t1niYUbb
Sf3E3+BnPw1vtkN4UP9T9+Xin/kwDCjsEiCeUAELnyc8jiF/PJMEmMTAx4CYjl6iMHrhi528LZo2
Ofj5FELvmNPo+Q9ZOhGwPmUEDrqVTinCeAlzF2fG9qAUaQFh9fGFw1Vn2243AcoKrK/vHGM0vRo+
SRVYczPjMmoNO3VlqTPi9dylvIC30Q+X6Hu2eQCcbOhX2BtHhxrzCfaEXZtsWN2iVkGX/Iwam3RU
7PRp8htVwcdPBdrER5AerGCkwG9uU/9jJq+aXjekwZzVWSab4SibOfaGriliHUQ9udCRMgFrQGji
bCRgufhsru/GsS/hoHyx6zKF9cWWwBWLqV9gMn2xC3Z6ndEj5C/ATL/xHVxDvZdks6N88evB/wGq
chtq149rN0R2liVniMqpx9juqXgm1njjebFdrbPRgGHC5VyBZ/cRATKjd0xq1wiCtoX1QFSx+G9p
dD+36gA1F7zaSJrUtXgcEKD02L5gfBusi6o7LzxQXUMFoTlBkxnAqfPrCKyQld3dOm/qW96n0k0v
DNJPbs6n9XqCkflC8Ytsxn3nyyWarHxPyxaauHgLeGXUdY4gS5RQYMlE+OU4Rl/M1+STjppFnl1L
EiJrfCi9oWg4cJb8q+BWJUrNJXwDX+KwxpINDSe8Rqa1w6d7dsoRFFwQxwrwZWW4qc716VioHDIx
MHYFfVfVwZVdJl8S0JMufJrhpAj+BPSk971+yfN8Ecb8J03eLn/zlaKcY1M6JgVfOcbd6DC0gBud
hCSMXfqqVGznDZSNV6J51A9KmR4an5pe6yrh8umchYDXeqCQYDnM9zhjkTvElhpcf+UKqQBf8KAt
nW6YMcVF2vxOK4ZAttcpt8NEx9ssrlPgJ9Yx6dh7mAXeWxOHBVLd4nwlRMEsDQkUpBHQ/e14vb68
cGR2r0+MCIzNRNy/tpOqKcByi4XmwsXhwmDIHm6wqkuicoT142IUW21h+m7xbQ0WOvaCqDpNscnd
duKLRjZ0BvdUOyQSULq6WOXVR4G6jpvNJslkzA79esq/fzWc59fUVvL8QSHWaJrPE33mfwMS3bvf
fI0yCG029o+WBfvZ479N+iwHRan9VdDpQu6crMan9SR8UVsNTxbRuoFUNvS+yXpmtT3SmED08q2F
qPjveDXIjiiQ++N7zOvVEIv6Zu1SohS/AB4Pufx6ma1+bRfNCCYlL6LdVZO6adAQnXCSzky0fiE2
xFmjbpy5o1jPfHVXhFTOBNULLfvexsw446f9R5ANWfTnht/naERymagYlWe/n87xw4EXEUW/7mqG
igwNG7dvCY7OAxBCUANN7/wiQssPyioV3dCi/LH0NVM0j7JN43MF/ikMGGwXHFvKmI1Xsmw8BvOG
AEmPWp2yR4AGE3YS5t84+KJbBVJZLwiyyA6WnlcIcx5gS/fBFp6BPrYya3BVCMxYaxRslfvm1Tch
ER0GblpUX8cj4suB8s0dT9lcnwKhU5Q1cLqoch9ahXBoc//Wt5r9ctNg2gY6iYbM3NyMEvf4qpC4
ww6pIrCowmmM1slc+VkBBxNKQ2PgDbZz5NiO7yEV2PXcdowG/KG9vLcxycheNS3vQmirrNS+8YK1
uofLHgghVrjUX3ha04zSgOp8rW+v8/0jEm3wNAFLxIWGc9A9ySOHtzCiR9bY7kDyPBy96jOPp3SM
IVS2ehhK0Ba2sELFbhcJQRQOwSbdNFdhDE+ASG+bstZtVD7ez49wj4WQjYRvcBI1ECDlyzXYzpOo
GqpUSPQaeViNlKSut/OILaxARVx9G3qz4YQ3Q+0kiOElRzsbY2J0EtXeQG1TUblksXJA9469xdQJ
bGBrrM9VnDZ1UbXs0AkEesEyAUNxU08Iq8xCbUnOUYDdKbinU8xoEYtZE6WaU/tCDFwf3ClSBLlg
TRZhWdV1ua38mSpjqOuEEeXzVGs7PteHG1073Pf0y0rzNJ4+cdFOb1wyAikkzN/8elX8w0HL04uJ
rt3jL9kn3YAw/gsBnl2XT/bYf48l4H1NrycTSlmTGZ9klCZkhJ7uFYiupReCOvWrq78QsDKqbE4T
3t+SPEjHtOY+ISzdTDBDLMqK7PSdKpJw/LhPuKd2FRvLA0eRXtxDoffhyDeIOrObdoSdSWPixjEi
ydOofOfD8pDLSQJ5pIxshNG+I5rrtPRNdt6tkH3+35tOrezPK1Mr3XPsP6aMzdP3ybTUW05UKPrT
lt8w2j+oFO/ZZeMiSIZvMedEKgI3gHnJ3BzMpcjBv7k2+RYKDc7fWq9ksRhaYgpD7vEOuUecfGX8
qgTXy9rneObK/DNYSAi849G44YHRiBPpUFDFqVBbFXylPw0MrZ/OjahnS0IWWeAZRWjLvGEWW2Y4
Hg1xsqn+vXs5dloEFC+oSaysD+uDLcSiG73B8ELHsQ9jtu3bNazDYiRChdk4IxBw1/shTnB3w5Hd
sH7ZOfwKM26of/OxX02N8qhDYYaPMug+icUlNRqDIG4eAWjY39++4giWi2ilzTT3tb8W3c7K/X21
XMRdLKjZ83DO0TcNADk04dbNabByASq+/kqVOT824eenTtENm8o23DiFwrDJgOxpfvnSYg9L4n2i
Jll1njyKWkzgFSlKgfCstoz04xc4fxpvG49IajNHpOmgp0o9YJ5Hl/zjt48lK3f64k5gWK6QXIv5
6RlqsGhxVxd6eIMbjphPP+6l/Vkdrq8jTx5JyVS3C0+b2zG4dQ3NRGXblmIM1UaqrRrSBy9nwMdH
glk3rDsw0xL59AkdkhZrtDBA/AJah4Sq22parrNfkr8Y8oM4VNYEcRrzeZqzcEX5gILgHTrEafKb
iVFM1EDo5hWqSu+BzHHwvHGwjpWbRkDOZw5JhtSrFOV0Xl3oV2UH/XDWeXtgUIQQiSMlJr+WWKm7
cf9qYn0CEhxJ9/Kt2hSfORmCOQnYi8qeI158XTfpNAgLDmbN0q+onJaO4HpZb+B/l6xp8MMDUKTI
sCJjAyr0snfJHGg3JheSKoJICceKhLt2fINjcMP5uyk6HfftioBAdCuJGLC+JdKrIUV9wqSIF/ti
Ho4paqZiiJ23JVLXsqA3xXjrJdN1Jm2Nv5Ha15d2DRf2rwSgkxxn/AZVeD3hDw4MXyn40x/VJtA1
h2CaUaGko0CAF8cDSpSktcR8mAjXIu16+kt6K/izahDK661BWy2cssQ6Hp9dhxlx8rzvLGag7eWx
SglxZGY5SDEY1FFMfIB1HcazSImG3UlUwSgUKcs377R+f+wcEJ4tVqYNeHCOBDeM7swiJgTrK0If
Jc4yBx8lcSXYLrA6+ABJgJobR7TxGMnT6ArQHyBbnu9+Lr/efFhwmLtKCM56klBFwjU1F+sN9D5f
fYhkxhOtQ1ibwvXtZR56X4fkZ/8zNT6grPaWVM6DSTE4v5yCZ3snMGSejcd4Vpt35rrOQMsjL6ch
olQ/WPPYC09QB3Myqy6ofMJJvY39nSLyTeAmeFT7EGuNooiHKem7IbioH8hhLpg5ZaJevX6w0wUR
TlAePuQfO8KjwvkRyQWk5ut0dfnR6MeU4Yy4DTG7fJXHb+r2me+F5Lp9Lz8XYji+/ZONrBCv1ODD
Wotu8f2E1HFkjK4UMRPNh9xtxkmFdR1/cVXSkgIiY2IqoVsk4nb3p8EYbLME/7Qpsku08VyNE+qc
oKIUqSbzeId3KlYJsjAVELiREIIWsDi1sjtdYZdKLquQbWrmp5L6VA8qIsL7/DyZzHUYU4Eym3zi
qWm+I9uAk7tWKrVudQuXU9vUBMTCMoujets7jXOiPe//ErSWXT0wJOcQsjDK8LuYZKGGzdxK3Tys
e++tdMm8Ac7BPRTvueSENiJLrOfWVrQ+3ZNnnEIKjTK95GOBQdeJNJVBf177UUXxOCzu7o+2QPOT
8nw/jwDUbHP8YPkwXPgv+BNj/tah5N2OxigotfIN1jEnXTJiyCZIYLhzUrsb/J98NwKkWJCXpsVS
ng2auiFgfQf7ndEUaNNVZQRjwPrRVCv2HxSGdRdu3steghVjHR3zQD9BRakW1cfFObGtmUjcQh08
2Xd5vN5L61Yru3X3pfRwhp5MYS/fqW0RdYgWYBa3CAIjX+K86dz0VdmowlwNZWnpZ2dTSOMT1CCj
hfKwrXY2gnINxwfKxpFn/lTYp0b3Akd5oPgtLzUcG5SNAbe5mZ0Wvz+fDFoD+RoCqtsuwSFeMO2x
OvHFqo9dX25mNImgmYLfngHOc9/E60EjDh6vLfMbmxlq66lDq4CtZ2Gw2sIiJGHv4ZN6SgOXvoE5
Sc/cEEB30xDlq+aMmo+8RdyZw+jtJHkVaKjQ2JLI2cPF+z+4CZJ5PJuyCOrzIe1cyB8tpEV1pxwp
N+t2Yddl+aQcyyxvHOnlstP62bHlMz3P/wnIvfoZKLB5XiNK9T008/NzAhMqcW9ok0F881//pAUV
pFU34gQiobXb2HIiH1qyVr5xUwKs5qhXJBxElFECXXIK6GwZWIsCS5sza+QYEFUfr/1wKjt6dPWM
G8DFLk0hBMPFCfltMMtsgqQElkFi59Mqf5ckGvFQWJTFJePzNIem7G2AcfPE5LVaZ1PcqgpS+6Fp
pBeVRMcO1saVJDMd3Qysddwmw1nifP7zp9G2dLNRWCJL3vUTsYCtjxU+7wATm4LgGHD6zi0vjGNU
5CMILxYQhkb9lCAylcPXq23rz0BTEht8+UTuXy5DjmpKygaEvMR7VWpmu7u5KwYmOHx6BJztSNzD
zPoQJUaV2sg49d7vddd7Mz+lWRL0YSY8LTpFacmlTWuB6mYufsFQjbtcRJ7Z25umcn5K426hSFJE
I9AXZ98DuqVJtNbDjfiwE//H8gq29ecELNGJYXGNuzS0KIR3MVaJvK/S7mxbDTQNvbfEgF/7RzLl
D+dxmotUw/ByoqaUy8tkLigthxIdd1heeBWfJ5kN1EmP/4azgZJJ3NSItMSKw6i6PpQWK98ryFCN
dTjy3GGIyKHQobr/eFtvEru9Wq8OoTtHVCI2i1vNOelZdwh5cWfiRxIrh7FgbgqikoKnwN+NQIvY
a9nw2UNAd/GRyC/uzWPeWrmX+X8GdEB1/RDaiIyP0j/4dwof1aehhxfc5goPFl8opzrcVEO1sQfj
ZODZExEC4Ves9Sx9NcKj/lhF9WpXD5zwJcwzdIj2BSnbAhlgCV+TQ1ixMX9Hu/0PuwtjM9dVar8L
9XkxBUqd1T37aRaNidRHmZBYHXwC+eK3XOFUliKU9Dw5EcUNMUzsSgm94ThfK1d4HPLiiHT5ll+r
36kl3y/7Dfdt9l6UblXFcIs6SDDtt8RIe+Wdp34NsISAVA/1DyJtSIP3D+82yTgWJYSBgFXE9u3R
G6K+qPyi3vtL5x5YaIosbH/8ZeEhyWKEE/TzK+P+UWSYOi4lJk4j0vHDIjbmKnd5EZHAT2v/4Ty5
uACP5aE69MDSjmUQ48w3KsmDpffL8F9Wfj5DwnyrHdVfbcUo8UqpiCXgD5mXr02AldPRMOKtlQlG
AhST04dLxtkFZpXWgRM2QHwPgvaLb7bHc8EWONtibaEh/uUa5puzOHe9G8xqYoH4CTT262WA31T/
EDbukLEOL0PgIOnpnnKpB0aiCYosvvnS4gvJbF8tx0n58sUGLfg9vFvtapKUTNKWzm0MtVDugC4X
27rMvZMIf2BVlj6oplfbaXLWJrhFgdkZ6egTUvDetan6dJcpFJzEB5T9qye4yB77f77DabEJPnPH
Y5JrvLxUwz0xpiz+XvJOqWw205mlPykzfoM2CfpZKgt2ZDLeZwTL+MEqDo9h4ym+hP6M78BEwyXe
w1wzIcLAuapNxpAkLsrgAMN1zCDcrujwcNod7Hhv9Almrmb0yjOEEx5LQGNoQYG0pASrk4SHuExI
m8XPwxkvkER+wpsFyrPTMy5KZKb8W1gKyhomH5qYqExMbWJyURjig/Bf15CU6Q7EMlo/BWh9KZhO
V7IV7Ha/VeRkEntWkx/0MiOqzZWEoS8dbwD12hzbVnDesK9k9b2PSqnCZYK1dxUkPY7LD8dLxRN+
6JnIrIQOQbs3ylP6d4S3anwZM/H+IFtmg7IYBhh/JO2l825WbWkhthqmEdyPYM/1OLx/mzgRHc+K
IgxASjgEgAh81/NNs7Q+ihM7pm+tjnkbr65X7zdH/FdAqA6i0vrOMfaecwSY/yDKxshuEduk2Dj8
E8HdXEmmB9qFbl1GmyBgr+tnQ7af7gtR7CFnGsimVZfdws8BCVvtjkc6aAiTUjdl801u7ouNeDti
Tazkj5HUNNnqxFRMgKnuuo4doO+by2wKXdS1taOJlNbAufOIlIyH201GjOHIhZmtVfJoqm0Ri7HK
agLoGL0cOPxBP8JMhTm/Pb960obKp2ykzGSnWbLcUpLJSddXf91FrNbBRZTt0qMm2Xaypd3bM1Vq
iMJ9Urc3ezriGmNpcQJlgM/RgKwHAWigIzZMNycbXmD5Djy9//RXNUnBbr+iDsuf4KRW5uVjw6LF
TmKUUet4JqUo8A2zCCbyR/Fu+ERwzwuGAslcS9OwRyxYAiNhmGnEFWhM/U1fcVX5CTPDhrOBSJj6
0iAs8QRm5yiYjk8zB6N9rOQyXDinYRuiCgszXgnYQjJgB9dq7s3EIHoBzeYhaIQodsAX6g7uvzwt
t39D2YaqGp9OWWr7YThjAqPflSG8nGBbbgPrs08g/HY/1FxpMLyH+BPr/ToaH+8vHXxuEPJCEVbV
B0vs4t1Ciy7G4+HWtCjoFBuvm24vVfAe22kVskmKARdQOFmsb+ndJjqOE+ZxK2RfyMGrFgBCKHZN
hkhl8eRf8NRU503pGS2LpWtWy7WT1MJglAglhEHFMT+nf0e6XTe9DII/4ATQoVWPiSTg3G1HUlNv
dPIDkAHZINkTV1OEm3Uj4P45JmI0qHBRSqvGRK7YMs/0xZHU5/otjmt1vRVuRi/4AlLCCLVy6DBj
+dNg+ISs3Wt5IhUIVnNR1K4MY8ILs1+3z3mQooSrF4DgTAgHQu11AY8UPzveFKZlEn+/v/MJP4Bl
a/QHeQO5PQOcvsQ0X8B56c6T3O4jHECW4H6OUOqnbOzh0/GAPu9WXFTg6706rKYlIXHGnE4foR8e
hZ2ETwfYxUWLY7SnMwfwELpKC0XkYwFLwwZT5SJdU+wdt39u5Bgza2CN87UnLwov3MYWyAo4+xWy
695j9D/qohYkY7M5zEGecjQdG3dcCGdPsMVCbNQOgWSDMdLPvjXCFwWITfa7o7WzovKpfRdLo+C1
dSU03rLDbBF9xBIynPz8JnvQlhAgbi9wE+MuffiqxtQiEk5AUc1gWzr1AQiEAeJo+I0YWu2tJVAw
J7epJZ+nO1ZEu8nTNpZVOuPBgH6nuAyLusrT5PIOgTnf6sG+Mr4f11YhZ1TBgJpGf1lzcYdwupLr
opg/3Ub/QgLaYGfblpAPsUchzrg80PvG+0eEt+qcSk1c7sWT5Ez/7YpNUjbk+jEBWu+0cX+7XY3E
QDqfDxYbEr4VT3f4lvWYz+JCrh5Ys+SVrO2hknRXU5JDcHMdjLUKstOPI0iHl5g+w8jWx1olMqcy
qKI4CnEESXM9urL7x5PQjXm3xqzCAsQk/K4zLOeFkrO0TERoj548GRAEAO4DnyybrgPQ56B0wc+Z
3v8Ch6kc1DsJNst7YK4tL7iJ2gjdS9eilC1HPi+weRHhRtlctQUnWKV0NVS0Z1rEvMOc/5HAvBV8
b2hI7keH4ythQe5h3JSl7wZon8MThqpV/+LFY+Bp4eovKCmBQNa9Nag95Zx8ztva36nnQBEqApj4
HMu1aRNfwvWAKu0fZKs5NfWDIPxbLvh3IQIMqg0QKshE5uxPNuxUDOvfJpICEU/dQhOF3s+1BYoC
5E/ygfbUHnre/zNFBpf2OPhjZ3kvv38YAcraOvSLLYr+zy8tobrPqqqJpGYPE8BvSnnkIVJme0no
DDYJgWDe8SkqALqhl6RZZA7E8GUBUWdvVQX6v0kOtQgjoqIDAW6pfr/wlV8yO0/eRwvo5O3IHDoo
4JnxBOO59bmQHxhxA4nVox5Uxco7ppc/LUodj7lWCMqmbU2tUu1lfVEvD1nIsFj7yP38RA97/GQ+
h0Z4B5PE6Ux1A9TsWlcQu5J2sJaTXlSpkwhKBbmLZFCFwjjNONlh4kwQZ3MXdtfBXZszQJgzDEQk
B6TvFRIs4+5sEgD6m20jyfL8AdfKLifFnR3yKpaNyVb2qpC2JqFY3SPoQ6qwTPnXrLETegMQRCNg
u98IxOXmrdtNvkeTSV84Nv2Fk+WI6iT5oxulQhVg7aB9M1ThjIQt4WqYKCWCGRTZs2Cey7D5cOea
zoB5r3XoVKcwjndge0pACVZbCKaoBUbqHEQldNadT2F48OqRi0zzrfAHyLyb26MBC/CuWuiMKkUj
GBZq221MN1yWYDrNE/YeppTNKN56OLcz678AhFR6eNGAJcewAjZIFRmcnwgLI4F7f0uGJR3VBvzd
9s2iBCp5kySkZLfv9M5bLwNNFz8kz6MnVtJ/Yfb5KrAEXPH00P2DKKOROT/4Z2xLBpng0touzcGn
CBM+G0j8ddn3gco4QsrSnJumR3e1FMFYnjsI2cOnasDboIG3pIQW4ZOG9BDrHqTDEaQ499b6ppuk
DtsXtmP/bp+WnHc52YfvJKPjwHHG+sXRVJxjEAVk+AcKpEd8y+kJp/ue4mwIEydjmN6eT0/mL4LD
oDjOC6pKJfIJ5p2EUjS84IwTwI5MTvvdk/R++WydvszphD1Papw8e3asT/uEXOd0Mlr18FOzUuUp
FDajnpqpcXgVQ0+771c+W7M/eg2sD69JsoB9StPBjpIGzl1nokNpzx/Z8x811R6Vzu+VD+crtNjv
mEooS7oHvC8u/8fAyYg7b9fKeMEEOSbcAE3GQb9hqqM4qm+3cJ4csPFAapYJqhdDdC/QSJwzLp0m
rnIxCL2Zr0BTRM3X7Ziiygf0xKUViU2IysihIgs3Z1ExhLTtXx3pBbgzCyWMjXTMvRWjfADokxwK
s6/aE/YBYXWkjJsBhMLXlzQMQkpcp2zykAK99MlXyCFqtkmp6j96RkZLCD4zQWA71Y44ViIsSqOR
RpEzAvzmQslg8DmSwpsUgVe7LLqPQafZnO31rA5jh1HtHJ+whUz1zb8Hb6ufANbOnGuPjnOGPzIx
8XCGieMcEIL5/v9L7aMQdArUJXQaHB9LhdaEPnvoo59n5o+THAjU4GlI8IpubarBok9u/TF0mn0a
51s83OQoT8vplINoQheS+IkGDOHfQ1nkGncuGZcmq03Kf2utnLNga9QA7Y8Wl2w4pouJ3n1/Ieml
wjbYDq7AqqOwgyU//qBT9Z/WgDxpbsZ/HDQqjxLNpwvyaimMne7rknZx/2uxUUFodFrUZobavv8B
2mmnyOkoMkdXwxYNjaHohlNBQbFiWvUTzG5LMInnVZVwM+Z7NQCnSKEKoMfgWVD2WGP8v4ip96nz
8zkvkGuJ5KiY6xyGB6qydaWmWkl7iE8f9SPTBSNMKMKN/C/nlfQerZKdnugG33Rvjin5t6Ka1hHM
Bnk8e0UTH9Cd3eOq4JSDo3r58cJxYr8jUYYtDz7YV9GMAekIf3sOl4Pc1e33xachsvwNabt50lrN
38rXw3bhfAS+q4SXXpwCSFC6QyIQWA1b3KrdI2tZ9qRLaMSQlyLfKDjwtEF0n47E9p4uD9RIIT40
NvvQjGOptWBLq1d2CBJlyYj0RXLGKe5VDxKAIwhWrJviriiFTQWUageRoqB+vDOBaoF/D6hisIj2
z5Usnl9AvkHS2/sCIC+Zw7VBxHY6eifnFBd3Pgx6499tiFI6bqTkVkXZE8EThKfwnwyWpZDhzNoN
vbYr/5fTZaZphTlQC4Yl1WEde4X5+R306cGl8KIl7c49arXA3xGTA3iLvlbEViQBEKJgjoq+i4NN
yqjBUrGk6d6GumLfusVgaFGKsr0JRqVf36m41ozRRy/Tkx9QalVxViZ44QCicn6c2KH/cn5jg5k2
X7FH8L20rsbs4tWe71AGUK/hDZ3oE3TIudxSQGca7fTrku8l7/cxwyc7bBPpO5C69+FRmCek2XED
+5zj+cKhFUPynHc2wAwFyBvUuDUMtECG1+Q9hLlTBoxyKijoq5IVvQT0eyl9BZS5WMYj1oZQs+1L
4Xw8AIFd6HqFuZM09/fzkc5owZnjnqS0Pm4OWACdUp2Cnx9bo6YVLsrdMq8pSrO+1/a21a3tGQn8
BqE0vwNUg3Qwsj98LLTAt/qUeiMSJded9JVedT4wn9nfqNT6ecM6N15P4xe0WmZjN2GnHdwwhP9s
x8pPZIIA1P+8u06Z8QLmw8M4X6102YeK0FzXbfM9GQhZ163Y45cLk6Hwc9lCqDPFCT5xbycGBuAf
1UjZfu7g7mDFpEjdFz/midE0YTpo+0AFil7Drm/HsrHrr9tyFjchLqEIXk3cq5rJNT+VGWpn5aXV
LKwlaeeDDEGy0gY0qgT1StwqgNyPcQUkodB6qV7+ejc0RUmM3WdO9ObJhSd/2/9NtEaEcuGvcM60
pW9N4BRgSJn0MLb4B4i9KYoMr12PjFKE+W0L1f98zvOhkrxQtF9EsYbWfvNPGu/8FCOGhPCFlGQN
Bma/EQcaW72AgAqz/puFKQnIp2WZG7KGYmRl01Ps9wE1GN/ykzkD99HPZ60wFkS4/dcICsq/CTKB
UDsGhxFkdcDwxC2VmEWIkDvHy8F6DhWAPAThqPsW/gCPCD/5hCUE3gdAnDHCqAbE0xBiv+pSnpgh
88ErwwtKc36bQtRS6vCaHuF8gNZ3z0x81eZ8JTrA9cfI3KPlCEigKfSiHdK7pZ3LVk2O67HHDlLU
g1KUUscYZaNBbV/4RuF2TWDXMcMoT+p+nq+HH0ISvy32zkMYO5mMbiOkB0xbq0HhcoWyYftJZSnv
JFpEtaHDvuWYVCXbPomAj/tUsnQfBmDDWNf2FeDEPchs53JP8rCI2kKgG4UussnvLDPoiz9IcU6f
4KiukN2pLG6gKpnyIx4gvCjjvSzcc3RnqOcLD8M6j8NxgDxeOUOkb2d23h0c3ZwaqEYdqzort+Yy
ahTGgCChDpDkE09dTt+MYgi0jDu2nKRI/i8eoPCv5cSe9GKQzhzFNA7FePIOFqXqmQka1heD2unz
naAaq9iY7Q5LphVEi5xgTpt6fAGoeG8OpI90cmygdH1wPUDp7Ld8eI5aZ8X+QlzFjxyh3FkLfnq0
oRaOUvbCdh0loc1O1lc5hhBDSWS/+q6VO84udbsN5mxdFxTkGqA4YQ/ZY1AHK4sf1ymKiHgS+M6H
vH/QWYJOqm1jvYXPHkYoijS4vBdqMW+le3xkfSnMNTXCbzVgoKWvLyqzFsiF9yjC2fp/EkJTfSC3
BRoJuKDGo7hm2NuazmfqJ+yfAcpOo8Jv4ID2HiwlB7VAiX753g7MnHK9BvcSEUm0/fXp18jqAMTE
xNkIp5H4JkqRN7P44UCn49FeD0LEJ4c2YxEGxFhtLp1xML+r7Qys5kez0AmnyAaC6cd3qkqex/um
s0DCsCjxGmg29qBm1dGKjH2JjQnTXp4PzkbJlAba6P2n5ICbLZj5Dr+aa1Q+TaJw6yJBAprNbr+5
XmMZWaVKdk1iRQrxet5qtY2v1hj9civUwUCDCFXIrCmTMirxELCOCQ7KW8NqTlaWx7Blz7cs5Y/D
QBw5PaDNR1O0XDUZJP2YYMq0TBzPHGHazhiUxrtR60MivwFsJ9qOJ30X1rMnWGfKOSE6+COuLlnv
sxwsoBxjjhvCmdiv7THBvGrsBtiXti5kDTO+963ZCBS6z2wYGb9zAOi4sUUZrzvBs/8EX9qhQ7L3
dRREE2yFy+eUi5ig17IqQl3ZCPnt810GlASRT/EJBSLUgJB+Qpjx6GolBB0B2lO/M76KsVOzkwy7
DvwObpKbq9alNDab1twMR8OXOyDSxx+oJ1KZhLIVB+6tbMM0G2hA4tcQ+7cOw2NJIA3km6SDbC+L
M+Qu8yDAX2z8IIiYXJS2BiZzTOKRSsL4xvUYQtQEWp5cSp4h9C6OqR562IN80osXCvuOQQe3sTDT
0Fnzq5btqFPLChYwXdqd8rDkMf6St2iTTYwOKAZwwBuFSRuS3VIOHmVYnLav6yhZOkH6Zb86od9V
2EHVaoeTKyGMmbRbEb/4JKRo72XB3VfMmAP9gomBUoPvv5lawUmDc9TA9WH+GsKdrETiML+uGkdt
5TxpGSAFUagRYiLzsTNaFM0DCA1YghZ7ZD23B+7BlcYwt/pwVqXjRJMTFMgeo70m51pRCOOisb/J
2VwGtN0wPjIWwC5PavYfe7EF+d/pBB+N7VoI80eereHvt5LEyEjIZzBvYcXvhnqVizA1AcwjMnoy
Pp3oXybiSxx3qwlrm0W5fbPXnrMywloG9OjYGoq+XHEv29/lhS6PUuqPEByxUmrxc/+WvvgxIpNG
JxtXlWC6R3WGB+C/mcw00noGkQ7iIucuhbvffFqegAJAp6QOaZDHZIYBLyk86MpJi9d0PFFlRXWs
tnqggG8R5oUIwd+OZLCnFLW5ryvTPjLYpvZrKTi1fs6jGRgTeD86EJ8H2iS3aGUtrIPfaEn0G2jW
omKfQ2VnJoWQVWxrWa5lWcOxfvrU6Vs+T64wwPD4QQB413IlmfQ5jRfMPou1jcgDEosGRBQUbFXc
SzmAYdVmvpXn6gnO0HdMzJTtHVZdrdUQ0wBav0tN/EJA+NQE8R8vAJmrc/pdJVJvMDhgGs90vbbW
ItiPzUypLMJu3Nt6v+wi1eaCsSxLtG2IIPNmR1Qp72rsckTipXh5RgJfGYTiQ+G88lfbm+D7LkFO
JZJIpTK1V/RfCeEcVOE6YaO/HDZWRnhPDBkWtt2L2/u3gtMGm3vUMIl36LzBzS0k9HXXi43dtO8L
IrpVzVKZ2ijpSxLs/kbE85xZK7KC1oeKE5JlJFTUcm5xE3qTEwIqf2SnfujVhEeujRnub95CQVmN
Mk3y+nZkQPbtCQaN2DIuk18NBokcI5zuDustpLgRKLoJQ2WaL0uIz8D7AlryC2pbcdUy8eoR4c/f
sNnPMsiCMl2A3z+QJh0R29mHRSYvN6whA+YMNPCtVN68p31O1wVw2kHDceAbS5HqzzREaYItytpb
E/fxElHMnjAiRJt2m9C1a/fGhibG6/RZiWGzmg7q72UA8aekN5DHJMrDpDgwFF0Mr/ebaLueT/QN
nEYlvEtQQV+Q3rGoxGE5RZAHlSTwv4WIzMIGYhI1UYG5s+ncDP7t5rPmNxwqbRLx2jW1A83Cw2Ee
USU4nP1a5rgZHpb9wxeF50mV8rb+SbFjm/58WZXv2d2SQvI5B+eh1ugvKWo7MsiSEleRYTPbk86H
VJPjcVP3X6jAVHssJja4MfflDGOVNUifyspmkntWaldQ8zz/8bp5D5L/rc63VhlixOMS5Mdr5Sai
WnoShTuVq1yH6DNnUuPgnRJ6LS8Fi2EXeLoN/lpZeYeHRXIRkCAuYPSVt8sp77HTunkAh18y80k4
tg4kY2GNqDjQc5TkmbobxY0VSFRA3ARR0oZw1LMVbxuT0vL2xDUZ4uy2lJZxVEG6TTfRtSVc2+Of
zicirep0yUrhTntolXpQIC8s1re6s5U+X0Q+znygM5HGfYPF/MZgh5AV0kjyBROxqiw2YWHpLphA
I3UHQdHGAWarYiX6PKHudGIFmznxRwODasK2KeMpQBH96svZYUk+sZsqpdAHhdzH8ZaBv9cXwnLH
NyXAi0opregYxwBewEKrH6jzaVYnnK6ChuHQFGWeqYXf8j7o1xD//AlW/7bpmF7HIN7FbfsQWSHC
TM/U7+lDCTvG7j46T9IObr697YC9uG6LlW5b/lu8Zte37qwJGEoJPWWtOysiq3oaBwLd8AjVRkjZ
picrdhRcf57yQ/hDDE22c9dpfFjrSoh/v4D9otrZDV3lffUZE+fTkdojC6XErnAZJA8blirNkDbM
Mq5Xb5V+GBlNS5CQiQovvl7dD0QvnbnA7025JPzJBNWfTzfYYLEg80BFMP/1pNJ8V/Zhxed/TJRx
s8IKbRwpJj1jrVCZqVAEH2m/c4EgJcBDtT0Cb0LN4Tk3nWcY+PkYChXYppuiVFQXyyLYJpNEeWiV
5yDPHVIAXxykVPTEQnyWeeauO2t2vKTzTLoz1Rb0nf+Q/JfZqiEvNelUTv3QW1u6w/2FRXTnBJud
O9GEz8j2UfyZeGlWYfvpGZhKwTG5AlJYEb3bTMozHN2UmV0qUAEc5krIiLKoZokUst4qiCa1KOOQ
HHyU9jwKISJxj9W2xrvXN3ILFHhiz+NF0C3t0RSCK//j7ugE52qo8Y/52EZAcJFtUMLPTLnWV9Av
QO2NXvYUZRxq5cJk0tpNugR+yY9RICr9yISLjLM3SKJpTKCyFeS7VS929ejmhoHvcfTT2FCBE7VR
/VWnKBlNMlQg4DforT1OkFGbYSQUm33PUNfZsSWS8FykiHuLYx+iFkEjbxtxamEfdvT6WpoTWPaz
+aCJUlU7zZvz5fN3CM27cUFQeifqBsjBl73nG4o77WwGaC/2CQY8tNkJdrXjdz2OWCxvuxwdf9Xy
WgTOZFGnlCX32Yq6VHKz01UrIoAiQV9X8DMVfgSp5VaLoaH47om0pmmfuvE9aPNJ+CC3cJIBMACR
j06ANIk2j837+HNTs1T7dH8wXAxnd3mfFJxs3Bj1/ZWzb7JmYx+coooJmobC6BI+bd4v0eV7PS85
bDEISWnBTNeCzmc/AehiWvSMdGHkQvxFdpBJrdEgwmtH9OjAJUEG23AnC1W6B4gVWX3jwM8QoKmH
TF29tke++JT83Qg2qzhd8VmWy0A0iEXykU8aNROq9DyImCQPZijOchSLtryDa6weIuLuTKfmuynb
PxslZBtRnhZKx2IvZpHdE6tkbbBhMlksroZSIhIDYPSi5BmHLmLdlOyNIwlJRRtoIlNQSdTwKdrW
0wKRD5N5ilgfBjk9tORN0KrOnA2El5x1L8IWNxZF9cc3mPcfvnFYFWBHEO3L40weRJizNXWnggNj
U8w96JEbiC/oWa8ZheMWWctaF8kHfaztB6AHb1ZGSvTJMaEAmDG1BPjgtZ369od7Ctihx7Xh6BcF
12G0f9t37XynSW4vaAlwoWrt4jGvgGrrecNBELQe87xpnDX/dAq2YpT2+Yk7G83f6UT+XcReltzm
NDacHR3sY+su0Y7bz3hCTbMvmBxH2aF2Yh0e0DDnc0/bhiF8dmpqLnkT6WrF3cNds/7nWLrakX3m
r7/JSSyNcymi89EaUplVWNYUEl6oDvtTjKVoabPjvE4q7C8jn2xagtuK6v3KMppTqM4jl1OEsfSf
bQUO6MrgH9MAD3YN0lvOAbCbsWeMafVvGkukmzuuzpBLlpZLEyNLRd7hx+xvn2Xs6avKkZUf8kw7
PODnmwv+3A7LN4firarPtaJQrLSJTheE2qngz07zgnDfRB2nRe2wbtCUbwszihpP7ftC2Jw857sY
EQMjCtlXgJU7zkYzP24LORqPRCThBoY28loPBwJhrHkxdQg+Q4jKsD4XQUqHr+vLb/qIeKw2kyyV
LzkPay8XkHIRzCwUVaHsdZkhSUK5WjSWPjngfvLphf+0oE4DqGo4u4/WYKxP7FPOFbiAFKK7taPj
EAMuiidN8Ap+7yB8RF+GaPfzAHsXrm+IrMWqymFBzazx+vl3x2xlxG0UEdVSdkBdwVnBnho3fh+q
ym6Wrjo1uiPAV2uThvLCxeUuseuKtGs56ffTmq2mEi4fn+n3IbZjtcG0/rWVLVCCtafR+HaxNO+H
S2J4b830wgScxmRXRwCufvRlc+ggvAOiJsnHQTpoxXdUSO0kH+DY/3iy8ep41MBHndlT+bWJR0gQ
jc8/7bkUN17PzAWEXfxYMYkRvfSqaeC9xAibjs1+9PVWElaEtvpxRzgkkRsai5Rm1lDLxINto+Eg
Nuh2DBos7ulHU27rXTAVMMVswaseeaMMuiZ9Y6LSyQo0SSooxM2VqM6aQSX0MZUMBR2uEsKLS+7h
XoHPrMKMJD1tuN5NjAA5NAdo+lKNP78fwS4YBRLUQjFME8ataXQMMhIk6+BlmXhYaOuVoCDjpKiQ
/lMl1a8+lkehXgXC9yRCGQLTAXvema2vJoxtWj5Z5iJUdLmoDcwOoXc/36DJsiwJxeZ4gkenzOks
GBtxB8641HhOTFQWMA1TEof3EtiCv5kYt52FtCxxCBskPNMHk8gDwq8DZ7sI4Jgzcr3LFuiH+XS1
V0/D5g9FoyG3W1oA28AgqtrtnRYsvr7+N9dkLQ4HUdUtyWx7XURpoVMyHLo3vX7lmMYCzklRl7+A
oLlJGz57iMt+CPe1Z2VncvxKdkAv2pBgDUYgkD3yU2j2vTwTitjN9PgsltBVUtZLOBo6A4kiFkn+
KooovyYDSXH3+wAz4dt8UCuKoGEj/8BRgYTL4eJhuZO/NsRZfWlwPLZjb5eJMZl/byGSNojY5Onu
dJCVqGJCT5yLblI9NYbHw4TthLTxmI4ui/HA6njWB3/QkIUPBFYKjHM05dvOLGU0ON0Zg36UtIoU
Bx3wl6PMTKCLcbQBu4aXbMF0M7iEqEjbCruzf0RSUzoRAwCam+pFWgtNUCKPe6D0oGSjcT1o+0eQ
6yel9pw+N2aVYWo1dbTwXZyB+9QQU3Fh0ZRFI1hkhjQZMXT4Qj99HtZ22hZmHYQFdHnAuUFjQj53
lUwS/WL294Zual/aYdLf03GC53iGsjn0Qe45TL5ht3QJGgW33mA1DN1mWei/YutGiE+kK++X4vnn
MmoMM/o5tiqxsD+OqgGNfvUcbs8/vm9QuK9Xbcwzq2L4TTLEY9GWBhUZdkbFmLvrc/9atnJ4TSnU
4F+mn3WmuXpT29YaJODEA0ryiyKywslEPqRP+WVwxwSiF+1W0IFh/UcGQAFPAjyuqqEvfrf8SZpD
c2R5ZF0LEDB08BHtJHWqwonUahjLW+tIRmo0P4JiTmsw1USy8cquxTsqmsDgELPAwaHElQwEg4T3
ArB4uug/GF9nATZ/YYsR4ujnqkk7Adk1/LnLSSrq0Rt9FmsRny01hUOZF+WZ1wOdAxHK/Rn4WEIh
jbhNr1AwuMghYF5a4tnloLeiKhFyXt8UjypGB2O8da8NUDIz6am9SofmhiZNMCuWJELt91/vBgON
uDMTRaCuyI1XuTWITYZM/QMsUyksT1tqHnhfG8hWDs7qZzUQW2WKVOFX6VwOhwyMzvToWJdtfP0s
RvYKN+mC3OoRM+adhrwlc9fgUXEnTQfWgNC7hmMwie3VpLlwc/Qyi/qk+NOJnymKhHcXcRVCX5rR
Bj+8qmupFmoJEddluAopj0JAlIPqaT4Qz7SUf89cxSDfdsRw7RfE1Zfj6+spj5O4Mobu4L0T/Whn
fhQlS530bpIQfTaao6xqBoSF/yX4qy4IHObTmj8sdN0vJk+l05OSLDxioxTUawhJtrG4rCdwrRxm
OTbjoDY2UttA9Qll3H3xY0/+iUdFCyT0fIdoy5seSccWWAtI2cb9QbNC7ikaMi/j4VX+aSglhHuv
LDogob+WoZn3Cga64uv9YGRhmX75k9d/YCh1BMsCGY4s/YCYeKKt/bs+mRRKyXiXCpifyzick1Y5
QbCyROMMK4J/01X+PA14z7Stgc8qM29bcq8ORIerPJpgp1cO/d6Ddt3W1rRL18feBcT7sxKXDzl4
lE/IrCHcDnBSyKrGRIlYrI44TlMP3F26ZleWIvBXIkZIcM09+JjA1fotzADoaGG0PzZNRv4fjIcZ
XPcMt1V8mgPJIgKZj3AEdssOSmOKNOWUItZ3+jH5xme9lTbqC6g/jYiqYZXhFftjPHTx+YkqnRLJ
S7ThFils7/fHY2wjTRemwSRyf8r9DF/E0eJKDi+KTtUf3DpyJFyKOzBq6I92F0l7pCT0DnYN5qwW
Y0RB0bosDkyAkzepRIfGFwGDr0FqCuGk/JRpH1I1uyXVUXgxkjFD8vDUBqpWBZR1qwMgd+tQO+Do
3vt5fA3BuZwHHpYxeHsY9Ql0Cbqr57194Ywu/XuZXMi2fL2LmWJlN+UuIJ79h7S2OgZbi63p9rBd
kzs+Px/RbIwawWkbv9Vh/DpLHPbLQMj902dR83cU1h+2lrMnG7W2L1C7fDv1tTkRfuYz8Ow8kXs5
Bm6U2oPGTJWjJyrz0FvhWYrxFy6kqpAAy2jZhOUYmui8zo3LbWINJHiE+AbQE8nzeB9w6EkxfyXJ
4qEDFoECw23L/2dpuqfGFTPHZVMfItfZTNU0XOgjeEh8wDpnnD5UCchu+s029nqTFRsM6FSy5sFi
Jq1QGb/xAuJ6XvZhEvolT52pJjjCuft+ny9U8LR/rR4gENnQMhGJ6s5K5Xc56N82MvRn6SEzdYH2
HrLYcBflwK/5qLKMa+jfRv3KFMmISdggWck3zzZxF+3gmRlTNhJlGteY4cgkPQclF1y9m6xjz7Hj
R47XASqT/td91sNGXZwcTA1b0mC8TZVt4MZDeIKPD9oq60DN8FJwZATfmk3rGjTIagEqx4Aey9bY
ZLq2/KYE1yy++Fs2DBl1fxJFTNGH4lj3rZPs7KBLuUNXfeHc1kxBt+gpyWCZpanBH8ejRj393aMX
IRBBVkCyXEhMcO6AEMIhQuMjvxZQhlmDkxieXORD9R89mFDUdJiJ8hjTT+dhXxSuoZIIF1MiRZMI
fPs1Zmk+8aKuQJw8mMx9qaG3/7xFCBW5BHGOrSL6QQVPLE56tJbQ9Tl5JwsBXdi2iZlHpi9mWB5p
56a/UkaZttTFZz3R4M5nzEa78PyJB2SdFk3g08cPQSyw6nLdUO/yITMRTZKn4IvwCzOn/JIFo3X1
By2ScAlrhEoJxMMXo8Yj2p16afHSoBFlRczIOtXG+2zu8JmzhMMFK03jFjPicOq9xnRe25gP/n5S
itc38rMk2fWJuhgvbSAj9bEbZNVfV++hZu//0wVkHMkCEnNV8xGw6XgvBMsYhNaZLZuYuWPidE2D
prFsWZ0EbTa1NoAKc5ltG96XNlUTaWqrSjcQE7NfkxOlD10OsZmy2vPMvl3FDKXboks4UmDkD/zM
lJfIn+cFUc0P8A+iNSJygBDXtrUlCFvCjAM0C+EmYaLIFUblivIX7CHO0HqQXO2n0GuDb2pEr9Kl
bxlZ8nzCDQPohIKU0AtjeE+cJt4mfFiCXbDUav7myFO12A2lKMI7iDUdu5qORsSke2JMvOE8Pc+C
AU48iwRydeywzhjjy/M1Dr7hfkOwg64gPFF7zv6bywVOXblKC8nC4aD9lZiFEB5rbxusqx8ik+2B
hsSg4mMaAwRHpkVdCrKEbmeC0QpyQ1cNNVDcoRPHdMDIN+s3nxdOfNKkI9ZbriJiPfkxBVEf2EwN
hLiDeYpIyKCyFQVLU+2y4+DYl8REMMQdTj79m/O3tZW6+LJAzGXWAyJgVzOmf1imqsG7veMeMnM3
5vHAnhNLL2jae11yufelw4j1AzmAOPAMDhtrsGHtUkTopcFFPCxhF7Oq5ugy7ih/Fvm+ltbaHt4h
Gwh9inv/tryN0krxqi5Sg4fCO8hR5oQPFDcH+LJVWaBVeXNYihHt8ICU8eFRBywEQ3yC0oAOgEjT
Y2GfBKIXW5WOytD2+88gKHSN/lmeskThFUToPPxdjjTQU5goMXF4HTIj1hdeIKAfhLHtSR7ir7ZB
qAzJ767Z+Fo52gRMs1hsYUkRmzHEUlNDgkXebeFFzQj6QMiRL/lgB/t8RGB/v1b2P4py3H5C9LGd
OvB1nSFcIOsyMTGNE8lZLnbCHnh8LsSr8sohryEW4nPEEHb7amyld1tid1zCCtNoDzkzTlhrRRGf
pTBUn3H4oZ424OVUq4t7C2qciVAKYNCAvQ5VpOnLoCtdtww1DPJEMe+L6K9E+/a8y6BNuWYpOVzX
Qonu/lzhUOwA906Et5/mJB1JhuPVy2B2hyLB0q1mKFZgcWr7Ax49JcYaKtumdpycgD2Z8LdUV7Ff
sbI8Z3K58qW4suglNqVBYKKaHQdOyPY8INwtmyfhLdVD2jGNyNtq6Ijd3A0EoQhz+LAubaeq+SMk
ZKxpg4OYVdtPmAIQ9s9NWHVgNNd22PGxOlDWIgR25GeFKWoEw9AobqxU7BnSt/gPMAihO78ktCOy
NY+DF/AIgd7jJgii3abX7ni9NL7hoTJ/9TGOSF2vaA48yO1E8M9Krrqr7jE/hrFjGVyqX4yYlfFw
8rBLsvGheZ09Atgb70uDRuXYh1SRx/D1frR4tj7AAumuCsQI4NI9qjJ87hU+wRM0heubJyOFCGis
aroGwL4WlWaYqS9+W+C1Qoz++94eXWRKw/7rxpCZTh3CIhsiCgPVcJhRa70+3A9yIILgZYkr8sO9
EzMOZzOJdapx1f5B0odCT39C3yEZIK6w9kyqhTCc1bDl+EHoIudCLzpH5jTe6dY+zvFJ1KxXHd2S
X4FgVh0pTIXI/6epeO0NYQbAh5SpC75bmapAoOUlZz9cCsu29ZmgwAWJwrGc6kGisstE1dT6ZpAl
KjVAuc9/0msKOsLSo/dOrRPOfEul10Eje3/kT93DJ1zOYtC0hgtyul2pTaleMxILgU/f8UIWVfAf
A28M/cMwmEa0qyupGT9XKkCRp6eRxjiv3DTLmT9k/K+czJhrKvlg7nmhwcTAexbDQiRY9WI2Z41/
YLPdF5L1hAxMza/xqPQBd3IY0g2pJd/uvZqWFnCAGDqDF173t/mIFYfyb0W0n/hOfJFQavB0LrGl
zpPAi+YwO01J2LiBMHvTaFd0ZQRjSO4GgOeYWMfLVGO6EjX/GAe4EGsTozNi9CBqXrZAOdHbQ2wP
Gptnyr6XvkDLYFyJkf/+IZ+/bt9AQFWBFB+8O8s+MUvyQKnq37quE8zDfrACjqyWK7SNJamtuJXy
KDve48S8WRELxwMhxv/sLbEJ45ggxLLQTUr2rIgEObMt2Abx/o1JCJlIgpINzkJUbaiN3cqQ1J0v
XEuvsCgYpb8ymiIctvQoWuyn6mlxNpYQha8eZ0PfqAHi9ecp1lScrAH/pt2SfeTUddAn4cydDVPr
/xrBa0aUcE3NaIhbRgcVKoCG9Pf2g/cFfX3BhtzT0LqontJYG5bT/YMocz8DQLkV0tLQPLNceoOG
Xia0moKJfxoCkghb7y+Pp+QXNxtxJ7f5f5pmfcRPMTH3nHGHBcS7kG5XGawWpRQ5CVz6AD3F1GWP
3ZnOG22CW2dqIbmUnb21KJBg9DtzsLGJEfWY/VyYeKfhk+lneLCDmZx9SbyuDgIP3pzmYS1wRgiH
kbUvVhBSHnon8XRcK/A9Alrj/5ZJxKa6PYxU+CLnPLzLT2Pn/fZP6kheg2giciJTecgG0gA/pyYp
BKSQBK5XdSJFgovPszK5kybjOa5wUVNLCfHnMUsO62aY9cGi2UZlwPTJCkYDHdPAIO94I/JH6v/j
GYLh/GfboX9YuDks2P81hIf0ke3TqYxJynDnnHwfgg2ms/nxRkrqLEEfy+jC2lDQSmsnx0oMQ/et
JjIqIs+Lr5pvUfp8ld4+sbY5wW3zrEqEJI218qjm9fQeJs6l3S1Mp55O60SevPrYIvKa1Bt5azwo
6PwzGTHSW4KCzIwMfF4yVZexLuCPy7D+Tt4Tc6zKPlsUb7OF+EQ4zI+lmmaGxQNHPrfUDrOsYDSt
ym+OfvWWmTgZdRx3U3uYlSUcx0Yc2clhkSuOPfgglfoJIYsOm1x92SmaDBhJdRDn+izBcqIq+9uX
5911BulBsKfGe+I2KowsmpmB9BNeDIvlJguU8lmO0uSe5btgC5pRo08ZA5LrvrdNwWZ8UH/DRRgE
DCjpushknTw+6J+JTYbYSkstmem57ngV5/rI04VKVVbqDVKoS63/6Nqgn35MOGREaObIlU2Jn35F
ey2k+Ox6CeNEDHaagimcmGKaa3mnOKkmuCs2BNxhpvV+d+kfgFaNAOl8P3x/5d7YjIQBwQ0tW/Xg
7it9iW0hNcattnVSC55SWZvE1MV6dBChKBXnV29PbSYmRF+mQ3aVmj6x4e78S7uW0+JzaF3dlKD6
mmObmsAfQJS0qhOkdDcN0tzrLpK61+823v6+BqiJzk50xTpdBW/b3pS+J2NBU+6NNEJWKoVZc/Yb
gYLAkaRVmFsgqpt8BKPBd4oBXaUNtOebO6FN+wtp9iYXYPR84GRVUNgGYes1+rMVAvsYvacgHDvy
7zYTs1AYCPoy01HZcjOW5WER6EjjjF7Lb1cvr8+6ISBoY088DFxSujn+lc7rDYPzVts3tQMWxRNQ
AnhxyiwfQk+wy6bekW+2Cxu1Y3id5xngyZ23eyFseh3owUpjSJZ1KwKysLg3ovmddM9N6A1VeXHw
p6iiezzE3rUNHCqCg/BoH272QdC+r7ivxX35H2DcxVGH7pHag/KuQczMC8U1imMmCGVw8kjTh/c0
og5GHiqZh1DT6xcgRmhN4mxdk0UC6eupxyLjfz0jS3MdRq/AcTs/67/z71BSKQF184N8ebmx01NS
VrDZjjxRXUa2VKNvc+ZQhlFYjt/FiVdwIvuAzhTLKs7hoL0a3I+f8rZvTmEIfz10R4H9G3PqZWer
Q2E3r51ZT54mKHPohYRwv/VXIDQcCig8AyqV8QucZjZpJgCfShMKtfahYlcyTPD1hFKzzEgvqMGw
3dnIQkCtKEbl5kKwsb5MjefEoS6B08UoMecVnz9O9jnSXO2cL0MJb7c7Dm4vS6vyXbGrXo8wuGfl
pvzTH5elO7Kza7LohfIooKdFWdF7rQ+6bAPJS+dbft1MZNfbBWCcoZdiCcffwbKGzo/PmlNhRKQt
+4nY7id28jHkKQ6KW1Pd+kUFz/Pmo0NqNTgdqm8sm9y1s2w/0TWMKDqFI0BrFO1sSAM/EdShHEmj
ftZO6ttmXCfiUnqscidxfh8ff9MEiAF8+5tDX0kpedWjL5LS8wTySSu2El7m6fiHBd0XIYpc5ubZ
rXy5oF9hjFsgpkd4XIC1GqYm2uUoE9P/o+MKKgiPUcH/iDuF0mPQV4rE7hANiCpvT7E4UMLXpV3t
SEnbVv66Sd33fDxEfG9et8niwAf3N2Pp4i2B3IDEKDsyjBQ3rsruWLgfGc8hR7QQMCFPwVxxKyxB
gzakrJbYD9RZdLA/z+klSY6iHmrG7GAxFQd0/VzjV+rqPOVZ8if4XsgArhrGZuX/0HyEiNNfbW2D
U1tGJasmjwc6Fctp2aNzs+HzWxIl1VPbR2oAAtVM0gq5vFJ78w7YIVUYP0vEmDBUTaXZV2VyKsxr
krSx2LQqWm8mGo72pka+KLBAX+5cmT+h2LzVUF/hGkSpJsRoa7fzdeouV7Y/fFFn2dyvSLOuYd/9
pJTQGsvT8sWqbJuOAnDRvQpyZjLRt0cSjCENCnbuneRvTMmXjDsyUGlhbv1/83HIGEEcc7iuQF3X
G4l7Iod5KPWwXGjIk5LbVSxhET0L4rUKcy+CTPFhWyRdeZHxRIVjVHDu7UGfmyaIrsdbw6TxW0+F
0kQF05mdJfqVVxHLrEo4V61QozKsKeem+SIPUhDwZVcD0ESk9z5oIWjc8sc6RDWAqgIvI7oJUsEq
puJWM8FOYGYEwOgMLDvKSmob6Hi/rCBF/uRBRzWvvR2s3ixoZI+Cnls9o0EADQ7WNNcT0Z9BUlFY
tHaXxWyoYHwUNwxh00UlyzysX3WrHIvPa3yrG8c0MPT0MmFPi3o6GskML4r2DfyvzqcXIueVCpYI
PHCRIefjB0sPwLqDJJpFYKq+BS/ALhg1vnWwauckwCUNemWMwVRBfgvEiQB1yMFHbeEdY7Y8RWQr
5wfIU08W0Nactpds2rj8MJAFrEtftOOsWlijdC1u5u6910MjDnvqR3k8zv3D9U59flLcK8muAjKD
Ok9dHFq5omMBw0qQ+X61jbtx32GgeeV2bQlKzTVJC3LbrHdeBr5yB+yE8eV1rBkO22eiAavN6KWI
oZ8PmE+qsBNp8a89ZjmeH0iJiNfXZSp02jw7Fh4E+EwkIjgnEoWKS/JcotPiP1nzuzaTKqxNi4pN
QEhibN+QrS3RHtRO3TwgM0mGhk+hSNwk/V2SNSnv9U4ceVUa0ARYvgkZlJJJJfYXqmFqxexmIpdw
Ws/JFAX4Tq+Ic2bkyY5/JR08h//2MW3sv36qYclRzmRWE5boyeeDKu/dWMbjXZqDpOvoFbCB5zDK
Jd7YlTY4vVpL/Pr9LJGO8REw9b2bMu8UjqmJqPc0PNnXyZMhm8QBkqqRTMedzqilsQ+8Pp2iHIt9
5o2nSuHsLMXhQ3ooFoTh6guBEB/UZyRELoiIuC62szu45BN0CFxrMk5NQdGTrjrdQUIczxpB46Hw
lOfex3yEhsI5H5xb+VbvHFJr2HSvQCnv1GlPmbXyhSKR/JkhNG2Zczn84hRoOTJ+7vr+B4fzyf5w
MJm6d14Ohj/EJkv/fj2ReWXqttO14xVvKiK+r0IvlETMssAmRaKU+IUgiaiOEcqh0bRXQrgcbTBK
ASv9c1O/ff0MasO6xqYsQ5n7Gc3fH6ovvY3NoO51qr0DuBD7fzUiGGO7abmIEMRq8qCOBvZ0VeA2
0vVm2t4FnyqnOjcfXBMBQJNkBR2xrUCFaXCSDFZhg6QoieW3NOFe8LNjUHdx1gIDXNZb2Bq1Hf57
gs8+KEBkXVs95b7BQDCZnP9RiEh+RCOryjjzHxIECmkDyf4tKgqk5p0zHxu1j1ab++sPHqyT51cP
8XnfJVy86q8CmVsn6RMI2Eikhmuz8ingrc/mYPPXtqXsOrScvtKr0gK0wLlScxxAFtzwcDi/JRS9
MZC9p3AfpvywkeyDP0TKxsdoecrkJMBfrHGyUXH0BxyvE51pGmdNE8gfJO5nAsD5zOcfavl2zv/z
YXl0lwadL5qRbSLB5jRc/m2YpdBUloEPbxAu8QeiULeTDFQ3qJ8ko800JZoUOhxshfmyTXRjfqNA
vZv00rMcXAYNysv0Qii7AH/CjLKgkOEfMB3959jxHJ4P9WD52i7XB9AxP1e7wRBzf+MEcnOxTJ9M
B1SL3H8xXep3UbKF1toCCh50JQsarZabLaL+GHZRRJbhRpo8LjsKKKNO/3dDX+J8Z4SEWGKizUaA
X73Zr3B3G5LGrAuoFmao+R3TqvlNuGccphKvSQ+Grv2sAyITI8cX6aDXPLLVK63G2XbN7J7717Dp
IDX4rZgHFhpqpw7yVRbQItTkD84Z0PblUA1sWNup1SwIrpDT8k4QgMh1KdbsyMOOPL92EZdDwpMb
mr9rRCoyGj2CgcFRDytdyD1KCzEExTRTva6DSnjbuYC3eD5/daIbjoBdz8WrJ0B8HuYjcn8YCvTc
71skkw/gGjzdhikJp9c7sdvLjplukpo/uanB+V6NQimsAQRR70wgSv1aE5ueB9zYdLgMUQp6KUBy
C6fu94rxiuVgC1Oo2zE1HlpgJLOf+E5tqBoTn9w8+P7jqh7sopsOBWeT36jaZeiXR43ZW7gQltwz
bazNw3knHvD9FS2/+sZSCHbqzTN+R7D2MAlcY3oFaN61Fa8vehg90Jp3p+S9VyOJjrFOgnKayqcX
ibHds6L0k8vfX9CCQR7O2J9+Zo3VVXud58ecUgrlm3uprRKGyeFf1gNAeGinHw30XoDYAULwCQ+Z
ubjMq4OZ4EfkGF8IEltkTva9+vSXSm9yl/Y1KH1SnwVnqN+uDfmJOeZANKUAVw3hegM5+nGiIC0m
ZdecB+U0SD5miqMaWP4HZyWrGZYQk2cHJ95iiYOcbhSy+b+GcaOxxqpPrVr18zxKef/jKlgpa+q/
0p3QhE5UrJvfOzWyQE9cktgqGypBNttBTAzWldGi6z5GO7asYL/xUPAOJeXyEt/xHjrtd53EjZC5
Fn5XsgU6epZzFJPVqIBoB6DEhaBxrCzMrUYp5u46MMDO4dnHajCdLxZk8yFzvV6hzE/+F8o/c1BN
z4KmRBUSK5zdG/YvfHvEGvxIWj1a+W0EB2RLwGwuNDd0AmXxwaKjsTDOFJmpMea4qSO/H+/OqfRz
ReWztsQmhuzcYCnNYsqkcQDJ7qwqWANypmthWNP/Ka24qR3XOoPbm9bO6j40kZGf9hPwiRCOOpo/
jah9GFhyBrPBqku5g8o6G6hp/gvX6//CUvH1wp4XH+Mfy69LsAku3RFZVsni02k35tY0xV/ka0Dc
8Q3zyNgtCvUCp066mxeELJ60rrdSSv9hZPc8LCObvzR2Z/2N7bxQKLhl0cq3Op/o4KZbUqIOgzXw
7LakUPtUwngZPLzC94jp1XTK93wlmiDnY4BqC4wjRl5qIl/LQBvTZYfNQwQ6xi1yjpgeO9VP1iop
OIfY3mmdrRtqwqM6AUFI4xlWkzwAoVkbZc9l/3eVlYuyR49Tsf+D31UA2a2C+h5zkK0Md0pW9r4r
JiJWEadM6STcto3HLmCEr27qqjHd+RCVVEXe3tAHT+kOIxLDaP+7OuKCql/fjSv+h99IR2RlPGAN
F7Zs1IVtUOQH1cDGBicnr+FaCsAmOn3nQO4p4nrnjk4nysoZ14W7Vm8+bQK6ISAmHh37ibid47Y9
ALkqbTBEIq57lHBkomQjTxqjHxxmE/Nccllot/52869z33J/H/aGpRZTem/FcpxP2IQgUMjaO0NI
D1Nrbl5IPQ+gDjO+hf918M2kbqe449KNOYDgoXuDaI7viiG0FqGv7nFseva1UgcIM3Gsj8QuehIt
IUK/H9hPZIldtvcJB3yhTpX6dcY6b0d5dP2C/unzym0L0xQzlUYDvxlG5LiOAgKMpUlGdXeVYCKL
V8XVVDm3QrC3j4O6/vQ3sjEAo/KWrwyGzincjVebg7JzXGAFOwbtqfSrlcxQ8ccU9k13Gj4KyJTL
CyGe3GVBiylAFVKaBaDTYCw64xV3XzaPHu+zVoNOoT17loTq/qaiL13heQZBbDP14X5kARQKAhH7
UNJNuJ1LqZ/lpCr9PCaKEAfT77GtKAM/eBLwlugelr6R//LMUQMxxMLl/O8mDz+sWOwED+svSn1s
LL2djoEC+Jv2olfrpWxtf5b6uRje6fsmg1RUx54hyrF6sbj4yLvUdIDWu0OpRjFeloYAmyRFupN2
PTAWC9YhZi82HxFxG9xlUR8YYHuRl7X+c6sp68gu0fgRqB+ZNHtDDtb6bhenpmqvgOrdhIh0ZjZ+
WPvpzthpOkPXy3picmpYJXeoqWRzws9lGEjKG3w1Y/kSH8MR2JrxfL+6LDuY2AFKgD9ypbYrRuEj
ekSn5K4PdEQggYpfhScLMdMPZsp9GBNqPM9sk6gU8wIXxuBcxVosl1oDBLVY06Dfw4J26Ix/RWWy
oXomCqQXW/04d22t9vJhnJ38/J4G/bEJs5nIuokjVVM2KBuo3rx8wnHFIt3G79MLHieXkLc9nTwp
RqzAjqR3qqzVTV2eJP1qTVinddEIuab1+XnuOpmADgyPzU48ASmyQpuJbvVDXImvM2yeFClIeBaz
k67atVCrBmmZU2srx/ZrVb9Qa+MTGJ0waNQp7rwjRAlXFfFiZVc/DjW9Ij/xL0Stpfmlhw9RsL6I
alWtPtlnX4pTi25zPQeQR7f9H2EabAc8AYN3PEa/hHPcG+tN/MHH9Tph1mbGyxjo95MzlVIoqw+5
Gf0hp92dgmbIztjhl0O1oo8ktbip169m7Vp8bV6z7WSSqX+vBNrDUYtsOtOtZbDgZnIu9XrlPlqu
GUj7Ffeu8YeBGx09oE2iyqSMVe3NNsoIjvvR6cJ3taedmLVSeTgP6slWwcx9tfAselp3OMGg9UeM
KOSyXPFYSlPAH9lrJRYNYPQoTIJ6zvRglzPpDp88tmir9U5mThEJa+1BBvCQtZEhpkaEnESywp3i
f0rnceMFNo+rHiH8++5NtTXocAzuLxs6MA5EJ0KZO5k9L0l9V5Bc9vA84r5Q2dhL+1qmdfihEKnv
cu92LMPIEe1EMk3yrDYd+RGJpGmtHev7D89tzddi6LNpL7IQ9TQZW/i89JsmcIKlLqS19MuMt/JQ
q4FPtHyDugX7e786DfD+mzWv+TvIwyJZJJOYq3le+Pk6mC43NyhZR2uqn7n4sl/VzEHV5TBmODsF
NawjD0k5sgEFNk4MCoIW18mYyV3/3v0bLs0LA/DhpCjl3mhcqNNXssc/MzN84qMhZ/NwTP6JrTCW
32LwoMzxSUwI3iouyn7gbGKqDDELJbFYlq+gaN1aTgU2XRIJZIegazqgvjuC8K0rikEw49/ADbRQ
szMkr3U+ufPPIrck6S/WURCukjE0qvtL4BfidzMS9c3qahj02Lp36NmK/M74elgyIOwd2D+LFwSW
mvACp/z07KBgfDzZljsG+n5LQNJd8alniWegG+rtRCUtAXKbNzripaTu3iV63ZhExyl2aaeNCxqH
1QwFdohAYiBXEccfftNe0u2lHkN91ty6QaQfxKZvOGzh3kEiiVF62rWP5YaQYv9rPKmeXdMPrvsL
dpBATIKYZ8aEXGbuRb3CtnUrBdU4bRrDgYfALKjbLQej2DuLlQU3ckpID/H8X5Hwr9GHX7IMcetT
rKyzJdmlrkM8yPQVnEKFwltXXlTJ9fAVn9HTnz0md/goL98d7Bg5Q0jNc/o5wb8OrQ6F9MdMx/J7
8CSMRX/nWttJs1OKflWQwinbk7Hl7ugEwMZ7cRLSSpLLiIlSzcl2PO5VUgMrr7QEJzat53tQuBvX
vwo6eVlYw7tkbDjPwHWPzgpeiFTAqGgT21DyiEqPUYPfMlwtdIYqOYOHBfLMV9r9+Es8bnfAjqbR
fTc7yhAQw4TL8WEOO46zlIGj5+ywpvxLYZWEc4rV1IsZTMn/uyHlp+/NNzxfEUq/lUrMe0HzrAIG
ug0oE9LatqtcNsrCJ/kHYhPmLfRg+Ywtmj+UWFg0c58BEnJzQyr35xl0Z5F5JtIDVX9PtIDDtlQQ
ulVPfyLiNlWuDysSUQt2h24BYAjqV7/JjuXmr5OSuTuO840ahyD/x6xDlCXzkoC4dTdr2KNJH6Dj
8Jb/LkdzTahzD8ojgtiGcc4X4OTgb53F5kGsG2qHUdfh9Z1naboPqG/d9yklWjH0jcQQ3b7qV1Mp
o0136TOJs2eqOPTVSZV+/ZNxaSDQ2Z1fmnwl05UDgf28yXhXBs+dIh082yjg5P/7hJDcH8Mf5k6Q
L3/IcUmR2/tHL7vEyu9aGajAVV+AH2HxikVHriM4/HttASI/kOAu0HOfxnVYD4x5BNWUDksybscq
K3e1M+SFCoN/Dq/LEtQhatsycSkZ3l+Z6JNkmknV+gLBvDwfvo9NLwuH8s86HBBxRFkGvYx7thFM
AkuFFK/kDa79OWfztP1DOlTsb7PIcYJPzszMhif4uLmUaLpFKGPrarj3gvrpCZPYNZDyM5r/SXXQ
pwJS5+D36LXEdXOeVQR8EF/+mtnb2nivVBuVmuPVziTsMn4G3bBmiwX/ZS6ymzyvl7vUxDqkxZlJ
Xoio1Q/HWuEE2wLJHxY8n1YznluiVYl8UNnQpmmK3sjBWRav6Knfi+70D9y8F0XTwupI7Y67wgZr
K/yYTrRa1s3xHK73ndMy7anZrmPsknqDemu7ll0MvR/OQ72g4AyBCYjsw0Tzexr6sIXvbmnEaznX
G4G5gPXEbxG6SNm3jLEN4yBZ3af5qNGIBi9cvGbNZJRkmrr11PvjG8adqYAy6FlweDy6Yi5Z+NKS
595tNk45dZs7ydFDLL1e/g8gvWOH5Gn7a+Lys7o8i2/Tj0EtnwNR6D/2PqyBV+A7V6B4dU5XV3LX
5VXt9gyLNpwbhgdUVywBPlp8N9OgiyOtbtKMJoWy9EZgrAD/OrD4iT1kxazBZs7A2F40xJFJ3lUp
8yobUc+X83n3rC9owRHOc7WhgjfpMfMfDiu2Y87PdjUR4QpChoyuPiKNiOLRDGRzYEphuLn4tRbi
BZeb+V1s6ueaLsHM/3tnQmy/gWq1HBka+lnZA8iGpM9eBbP6gtQmRRy3Iq2rzQQyxEIHd9tFw3MO
/Yb8tzEjt8Y+4wh8lricOJyWd9GXX8iVqS4SypjRiLNV+A1TU3pVddM5/FJy61tcrhCwRlrqpKa3
2FeaE8HUm6n5rCrVlmkUes5echdPkwnrcg+ACZr9Xx4zseteJcuy9JS1PY2j0GlowPR+l0r9Btj2
kZV1/alkno/yGM2AW5caaVVT5XojFi+lnKB4la5tl9M6KRjYB+b85ua/yg3WLxqMswy0uRBdegjz
EsAPt9J37yYcnGJh+arhOYCgR4oM41JVL7wUpjUqwgexNlLuxhnqr6u1UiJFfBlos1/jnXHwFBUr
/vTc91PZspHJaXiy2t16fYu/h3XgVVtxrIBFH4j5T5R3COefiZ0VD4D7JK45kJA/U5KuYRsoYt1B
gtEcVbZqmm8blkCjjmuzlDpF7cSDeIW5irnnN58fcs+besGM6P7PcXwXoDE3rMx/Fzq/laSb0/ER
9xaH6y3HxPLnWSojzYe476Lu1i3sjeM22KyJJihZ98a+KvISpddsKJkIPKaX985fQ3YdILBeFclC
Rj1rIJDQLv6WOPPqdjz/aA45/aMN9yVMvRiPWjAVc89/YE0LzxWMMlur3DREWR+UaxBivA0te4P0
0jt7Tg/d0MfBHspGv9hllNbZuN8vE/c72esGOZjsFGIL8C1sHih63LwUGv3zJqH6VOsylZpuhiSN
WZBvRsFi+7Ec3WsOlMH//357Pcq4+oUM3KerbqwGIZ7T+KhSekRLs9iYteiRXYr0LqviGCVSrxgi
n9NiSfS26ggFMXeE7hAy0HVRNRkBIhg4s+TqHbGoj1mYb1moLm990lMVLLWzMSN7dWx/9htRqWbi
9Pz6333VquBSg7OUmxD9TOkKK9muiSL5UKcosKz3ZX6duz/I5O9Bek/64GT0npLcbcyhLbD8Ahsl
LawS6xWzkjMOJGjIjVrs9WV5+220G2lMxcOSeDA5mri3WntsTMryUzbGTUXv6bzT7Vr2csSVMr75
AdwY8EUyUINxZ8fA8G5VRTTUUwuxKToUYuMsbdkiGpzb9AXNj0a0tgDvfPTYuLGVOVKhGT+JDCD+
3pHokZRO7ROXFhRILUttGp1Kx7VCYNybgt2Rmfa5JpbPxlz3eTH2yjFK+GjQMIVp/3aR8DBB+8jJ
P+28sEciH/5NFIwUmM+wLx0WcB/1XFNZboCJRT3KcdhGXopjyxl9ffJn1Fc6+r/nw9dr2C8YPeYR
678MBRd7FmIDP3ZldGTBikO32BWzun1cd5xB8FARcAcLllYO7KDByVWm0I8+4qmVkeHC1mRhBnnG
Bq7a0fwrIK2ZHbdgmjqYBXMbLxSkUan5sh4FpGGXwujvKhbFeGRnYMPOdwEc/am0PYUR+DML2Z/I
Ef9/wWxqMSTS+DQPD+uj5czakVWKoDmh/fWYMpj4Zs2/oCBT5e9jIUMxdBoUUVSpBQ4oJLEZCrh2
1V18/hfjGVzu3IkcrayCP6gl9vmrfiYHrYhEMe4ZIuLqBa6REbOigBeH99cKbn7n/bM3pmo1yDVZ
78y+7jtc336fYcHPwO+39xLc72hiPNjNtmrokxVkQW5Q/01/QsN9cIZXvcN2dQIjQ981WDO2P06n
ZAURndlv2nscopBE/E1U7lr5Cr9YN9XPXfUdvbYQp/3ouA78IRPGnLCitnFNAKSZzjxn/JvhKthO
dDUjiSOZKUcRgeXhWC888daCNLGCcRakwAWG6vArJw1hw1mUuPwd1in20BdbgEVvx+RTo5nAPXcM
4vgjoHtVpuwTfPePTaFrtaExcxkBroSmTrwtLt/lf18tYWVkL5HsN2obLn0JLcpJSBk6eS58DClE
1wR8CBq/3rlFj+p9h3IXp5kW0PoXGm/B+aU/9OGuxJpwXJs0/yvdSKnkf8n4LqRr6PSSsijIM757
Fb3+Ojfj7Ps4gF0OPl3a341ANGI+B7FyqtW5UMAw8b0QMfWYzh4dqIy+HJyfiK5Q09IgUgQx0z3I
qJPtuhg0dsa3HtTeSuBxT4wJ+m1fqd54rA49PSGTMGfkSIVFM6NrKOFIJ0RDL0SDaJOLUyjFizAB
qkVScQSoylkJEDoDfsSBNR1LI43Fg0+Gm7ZfTuOaoI3Z3h28g0LN4z2/c7+kUL2Viik1579NIYEs
0zJ8Sr4NM6W+fdg+ccktxlrFRv4e2UfrBMkvgxcbjfeUDjuOb5dOz/1WqVE9LiUKt7FoXmDycoMs
TJAcsmpJf3PtmpnOcJ4GHBJOPpMFJAiE2BCf6+CBVK8fiaUXMl9H60i5xoHfLg1yocc23otOPktf
T19T6KM4MF0R6Rf0VV4W7WvqpQivEmoxzplxzLNJNGtqnPi2gP4PaLtgbeg03kDbCRlbUHSe4FwH
I+XCKjzgJ7nsTbSse4kQ64JGCSDvpqVQxQudDB2zZghMbcdtYiB0LNy1i8wT9GLH+0yycWGiTEMs
QudlUxU0zTVpXf6Nrr5AFHKlH6tpvdn2HnvRAwZIPlSY2CZJ7kQC/zVTWOc+NSVEw96PNSOseL44
ISUyeBQphHekg0cUe6jAFjsmD7buC4OY60MDDjG84D2qQq0nMth4YE2cq6L2O9Rs3npUBdklD0kZ
h4sRgNfZWx7YazizigfX38fnBxWdT+SsPVWyBwhgC0pPPetlanXVlYEzTuIxehE0f22gPALksOOl
l94xpdnnh91HT4iiNJlqvJTxca0TWnDBKDF543/h/8P7QOJ/NNwJy4nWi1gKhtWVxl9agZBkNYQt
asjt4a1FRWtCbgYNWssr3Wx6TI5R+ddny+Fr5EIituBoFifqE12F2iULikpgWLkkZkmbWQebzAAF
IKd4TcBPEvrLL0a26S6A45ajWEfGHqVqIckkAzdZi+HP8dmTZZtx4ljB1BPBejWHJpaDucPV+sxy
Vm1DEuwEXSfqzdsDLP2Rsd8jzW8oDIQb8h1+e2pF3ThR2gQtyvJ2zIdtUA8Bq7EZaCHAhNT4Trc7
kY+3WooiDPDDC658huDjNGlnOqKAttRa6QnXJCXtO9kwkC1+6Huojc5URb/Q13ubFlDEezCcPwyG
gYzcPPLNyNrtepJ1znBiQUq2QnkGoHfv/452TAprwNHE+Dqp3XbFEAqrZ1fhdF9X7Mw0oppK5HrD
ZZHq3kXRj6acXhrqLxshXj+HGSNCkUiOhalCSU4P0eI9AW6io8thdGvCCLi5dS7Tl/jWy+pfn6q+
S3PiH8dvlO3mRw4eL5kC0LXwcKWxw5aCf/NXwdNFNavYaXTWhB9ZvZkUFzNGoUTfpblmmQ8iOCb5
RnYiPLySX+PTsAW2t2ogkOTPpxz0cvmcowEB+UImKGhf513EFedJ3Fs09ubh+hUL4LODsBYVENQh
jSNxHeuavrNf3pBcNnFAVqoIcQywXkHwRCIlNGd+qu0dt2Jn/EF/rmcQo1EGug6uy2Gc8EicNQWG
yjRtn6ddMzMlRy+ttqPZo7jlidnuLjPfJxAPLgYDMuj5y3aZQR2xcXXaukLYK7RiMzFcWhbhIqxg
Ov1uqLnsfU1cxIdF33Uio0E1S/kQ2fbXdhj7eKaE6ypQ1QPyN4yWHAHQuv/oeA9bfpbZuDRBo2XP
KR+mJbQo1cj6ZQbxGrlfN0vWTi0iGF4QALFfVry9yWzqmu+R3OJeYvdTsw2PQc431ygXvKjgFRIy
KemtIYFdYJfUFmrzfTkKUe0OYWzdvOFQuhX3Z/GvkowY/fI+0DF1t5q462TccdjoBQFPAFc/Tqgi
LGytsq613c+lix9Bq27SfD/JcfgyQ1s4W7+ItFZyrrNtxUySLfZ99+udhklK0HrssnFBy4GxYiPO
Pwhb771IAlWroZWupOHAI18wQ4FDSzrJUbwUs1KiPAqHjTmHE3div+tA2eYY0cjpdvSJS5gjPseu
OjWIMFZTYsLk0ZS7UfK0R+PhybDuJzmUkLX6KMnR0GqYmuK/1HtYULzAbdijCJe43H02gXFEdXD5
vHE5JtlIefVETHHFa2WHP/WF4WZj1IavPW1jR7BJkVdfo6TIiswXJRbZRp5fWeAGDszpLRRkb0gh
iR+aKTT60ntrVCTnpNfq5BHBGtsMETjkK40dzDhVueK27owi2EEVtpFlMAMyZRssz7ckjGHbwWvl
82+WmbD/5wCs+rsfnvyrB76UNonsf1qoK9pqQBYmjgwAJwiz5MKIYEmd2LuYH7IDRdCASMHk3Fgj
9mBiI/pFonzntKCJ4ux6S2HpOsG86sokJnAagpb6WSOrjBKxydB3dekY/CSCh0JKOQwoo5vUfqQi
1h7yNJbmoqhYdkS2qTXvrAX3SUyN670CtCMzD1ElFnRkNsXEsjUaMMZ5StKl3P/vmwJkn2tkufsf
oHQJqI6A1U6I9qv4m64RCScfuav26df8n7m9HY9LRQsKbhDJEYKMqI1r+8Sn3GqeqoRduSXNpUy+
8xBzBD4ZtBgyQK19Ca4KZJKYMdAKY6/7sXi2uI8qS9haCRjJMEtBEVhINdLp2N7LQ/Y9xwuxFdjD
W/PU5YVKKCkmn/LZ5vBDWYX6ynEfAuL0o+V4r4EvRg8VWuDQx7dNoQe9zZKEao05mpgwL/56zfVQ
Ttuy0iIQ/qUeQwkLUnkffzJwJU78Nx3zOewTgqPkZyxXcURqNZK/v94E95JQmtvUPtTjz251ohMz
0n+ZJK0rO6S0L6oGKMHSuen/6SDTwAtO3w6E5zifNkQ1CFin7oSVAJzTmvFH09k9wmTDL2tWA5Vh
21v2lAbCUylR71hXM0KPlKekC+KxRpMXKEB8VPA4MVkmgHtk17dqJK4f6SzGzfKOzc82bPLqLkQA
BdKwp6zgy49N3uUAYJedPN1EEHWFwufS81v3OScZBM2IOwaz67SZtTVk/xgC2tQ1ZwnBGs3ClB/E
DRibg0qr3Th3UX2dogU38J5xMslf4yy3+DXUD8orgZXcsBT4ddbeVQq0onN84bcPiFYAZxxiQP1E
ZePbUqJKxQS2y45ZsEzRWCbbcB/UgBhCjsgtrZNZEjsLjqCgir8SrabxbIrNn3oy1TbAL9LZhAe1
FTWcp/pRHzAdoI7WcHGyyZrplzqGkuvaXvg1Kv+9mX5brp/3lic2tF5bwLb2g6pjVCUxxhjOrU7O
mkY41qiEVnZNyiRBpYmHmbLWeNyVRAVWwSZUU8kPHh9U/vtTdwD2yGDt5JFzcsqxfora2oi8H06J
Omw5fJiJK7DJWuIzG/SlDbk35Lv/tBLxsQbIn8A2mdzTbosPe9Rsy7m4aI+PyvmI4/j4X9n3c0ol
mZiRtxQG6siQ7xbVredbAjULsVRQsk/Otsww3zxn6rjgV94D0aqzsjZ4qlVtMJEWP6ZSlL68OMcA
bSCrzxWWWDDgj3/NgGs5OnfKhsko8PEo5yHEttc7X5lX5k9mktaFTOIFhE+2sMzpQWcvXR1KLQIA
yZzIOhla4e40qwK8f4kMkgV6UiJBjkr+d/SIR5+u0wQDV+/D0c2O285KWaHUxeuzQmGjkOgK5Ghr
A3oYcMCqpT87jhmofLx9LDK+JbhoavudyDPdaDlAUWsVN3QSo3JLax2tpkCNGFrbhDHFoaSYFr6J
UTskDHeWObOmZ0C/ZDZRvjnAXfwjswm9w9BOFSNPfEPGih4M+QTyYSqihorKsvqrJHHu1PEQM11a
IyVGLqgK8XoU4zswGrTBQwiZ+TgjKy4uvklPu+iM3YhfH1x0BYNZaZvuEcfeKJa0wgWbTxJdKoQV
MhHe+jwq/6YRxACN8X5Z+DApCfiaN6U+sKDZs4AlKkzn1M0IWpTycmCk6QRpuzbjBdGaOl+MKQA/
U2iLnc2O1GU7kZFY3LP0MNAD/MjmpXIqmtM3c6FMvr0s3PJmOkdhXAFF1ZN1jlsmzQ8Royz2asPF
q/7XJK74iqV5iwGmQ5mUmXEUAGXkt3MOt35UwpIvnI53EJYhEzO1BXiMtxkz1uu63Cvak6Rcpsys
Dmz551t4XDD1v3I/iA4jIFVMTVVRGb7pOYf9+4N3Ml4urddUE8x4M5wvO4mgjAZLCA0q7yBeYnz/
W+hHhIqa5H3GRH9Eex8S9XB4raQdFBPmWVKFNgVmL5bQO6/9s+KnTIbb8Jj+CEfd/jJ6pwuwTrh+
sxiifk00I47FGhFL/GlSst6tkm87o+dePZoJeQOSYBkCQkyz9hzMdhIdRYscNMkEqfi2A9ALu5uW
JCmhoUf+WR6bQt6oaM7yFd5yLogOgY12eyjQVyCRjjX4SdD3ZdfsWaUz/NU0ITwV3ZQj7aLu4suo
W1rTs/CPqq4xnBK2zwTtGPuRj3PB9FEjGp455/NQK3yo5dn2TR8Qyud2IZdNmeWiYJpFc3JpU8tH
zrvqvcl3sidb7SQn+JOHWbsK7OHjuZGicqha+3gSKbRHwfHZJf5CQ4iKu0PeaeVpwDvR0z+LTFP3
jiopdav4jUy7kKJwPd/dKxDDA/JOGpcTBr7Lm7LMmRX1o4RYYH9PucmbHuuzkgNrDxHZDahCwrwg
AkAP9lpCHFsT/jMnJKekv8jenHNJgatb9f6QcjlrhH7V3NEtaJ2HLfwwtLfyNEw4q4l/VqbwTg3+
C3wRGaARb5kxxCETygckYTBdwRrlS40BdlH1B8mM8osxNys23o2ej8DyxD6mkVvaWN7wWbbugD4L
/u/O6Gg5SpYo+cDCTW7P9fYUHZ1LxxLwUqeTKIixen6K5bSHADybiq2TVhDi5aZTF+rRZMq1JNnX
O28kNkZMIJ6fzsUePYbSD5pfoSp2MgS7ACtSupAABq3F5qpXRPagUAIn/tDpiUYTMU7W0GGPkdX4
piJEsBtPiLQGnvPPe5D95Ne5lw9tvTqeMmSpE2a5b8GtFQR4Nhm3lDt/Q6EVpCe/v19bnSA13f15
0VeQbAlO//eZmMKZcWJ/nU+2Nuu377b3kguZOKIsZ4cKkouvR/DQ/eD47BNOJr8xrVW0Jd0isCXF
6J+VLHqOIrqG1+2HdEeZ5+6gvGW8vuzxEYdM+Ey9RRMNmelG+08UKu3wmmn/bCrP2RXjVqHut81+
KPkw3cdm+lFYYDy5vqyhsmwzZuFeTDUsHgfKAyhI0brBQxi91Q/R8c4PJLQDNm0UpL/y25BsN3XP
kN1sliOGYRlQjnERVF2t3rVtFOgMgicqrhfzk5nLn9BZe3yfisNdyqcRPjivCtfDk9OVPrabWHQO
oWFGAz/SkiWyqST9Ir8PJcKz2UQ+o1y4UOpBCw9/+6HuwvFCt904VES1buBMa779g/GSnJjUukvq
pgUTReUO5hGuNB5bygTMgaXDawCUYKHDJe0+qV7mN5y7ERIz+SwP6pNhm54/6M1yv3bFmp1ND5IC
Y9AKRLLxZTRyDrKb3idZhkYMmwNQDBW4/kBqZ3Jp9PdXJ+HbxYUFaMkBrZHtOBdUKb0HkUgY4Q9c
H4KEiK/3IB2yZicSGbti8v2SUb05IFb60I+wO1vu4Ksfe9R3Xco88GYVqfQ6JbPLtItYlTMLg7Sk
/EltoyE3H3FZLLLjuah19tsawU3h+BR+G6ktWNilS7wKjiZVD6mUZA2XBkeGlfRG6WrHQB87aLO1
Ocb91XpveWZhKeYH4Xp8M98SDf+xpJawTTmOIj0KOYigmKEBB/3cEfCTEo2/9y4Ixzc7RI+89aAl
g5yT9wsJDU576KZceviGz2vlcq5NA0aVWs+1TGlPsPRbAq7BtSSKspwCgxcumUd2w31X9Gj5oFT4
BAQe1r3wc9AJRD6orqoz4T25rdNejJm7gsuhrDwg9Cl89AHI0c8WrnsqqvbKwpaobwW69npjuJts
1qBgFv0tIUxq+6sL5qk7QPaiYM6L6PxtidutYyzccUsa9l3AdvW6wWDHIWV8V4WE9LMk78XsGdk1
uWojXbo/OdRTtjRsE4+7I2Wur7Ttr/50Z45f78uJl6orjz6veiDiFqBHvC2BoSwUfJaHZVIeJvQp
/ec2dXHKknDZQlqqK4qS1Q90t0PYHoxrst/4s6ZuozyaIFr8sC4Nh46PZgvnl6+UQPyIBRjT1nRK
56UsrUwo3aFDmOLsBriEEf8tZLc2zpsP/qZjrXfqQ6PrgyjGLXsKjbRJmOcrUjvMxHkkzKpyaK6Y
n0eNTks9sE/Czth2J00d2bHRRv5bIootD3BGDtVzqroM38ksTdi/GNAdvHxZwIXRw4rsdCx2nROU
IfZWbR7sjBA7AgH6LnMM5VpH85AsPo9TefB5FE5B+EH/xfy4QVAkN6GN8ArQrJtrOsAizTWa0FdE
xrAcD3lncN8aXoIMulR1wRWNhIIJKxUwmg9WFQDBRGtFUZ3lOGVMVgqOioHpQrfvParghtI3EIn/
GR6TmEkriGXY7MoJbuctbY2/dGjuytYCU5JDsTqz8DVd6MiI5151fmstt73YptguYDeoZ/uYPcmd
+tT/TlhHRwkxbHrnCWjjr3+dGO4gilVf8mhFpkTq9ndpTgAUS9aB6CtHtcAKajWdOJ4GOA3Kkg/D
962jQTpzyj6NV1BdBZlBeq25HSf8PSaRN05z4H3lZ0dlgJkRGC4QclO4rD8LTSk4YwwzL46T05fj
mNlr3gDn8WWyXtMTfeCW85Z0jxwFjveHDt3mpAPI+eI/h12ZkruMWhdEdDlazbOJZA17G0qQBGx4
ihXWe0bAyI5YNGIbSPiA3XoC2vebuQh2igXEkKMKwquF4NXJqHRjxgIEmygq0KlJUrsriovd0YPS
hgQa5TMXF85o81C4gWCSY9/SRDr1AzRAQzXUN2JGK1Gkq6N4iHURDhVtEKIR8JD0qDNhkuKkxzkh
CzmqBKILZjNfRnbseJei925b8uJbL+yAykJhTF81ycRXaMxITHEuX34I2b0T54pFD01sEsL/dFHh
G+FpOFR2CmNdXqOVIQ3yNmDl2eKX2tK4bUmbqNgNd6E2Zc+f4O2wZGfFOmPtg+/v8E5OaMUX5/W3
G2m4Q/2ZICMuWA26hSqTTFxUGjKhd+D0lG6oKTT3Ir8e2hX/glvaZSitsG9+BMwbNpRdtXyou3/F
NMovUNgWC71jtJJYtcy1eDPrFwzgaKWzuWPif+ePOoUvrquuDBvV/y9rWFPSbImO6o0touvQN0D/
FPyQGGOzomfLJja+c3i53JbSPc4q+YLqF1I1UH/PdGTIQ/ispjc8L54YeFjvQlz39r+1JW96fsWC
QZrPnx5a3bDlN1lQzOE2CO8u4faJPfRQAuepcjrcZWl63nLjkNOIv1DK22gCrq9ZSoU5csTjhPrB
5xI+wbxXduzmulFVVgKlQAs6mBaSEG3tXyh/PXy6MGrOhuvxFG8iJEZxmn4qpO+nZwI7FypNl68y
PNGjFVT8+otha5rLyT51rrjOhkmqv0uD4oXKqvQUDq/AUMCVGxy/DhGGsM1S4RT6EUiyF3jNc5D6
cRVAeMloWmiEi/i8Y2KEOFmBFMJ1KwLDZDOFWcg08udmgpXbxochnxzqionjNmrsXXlCjzJTnFAx
8cYNXnIPaVOIFJMXrwQZoafRNm7Qa0VVuFYJoCrMTjJVy9gcSN+1+GJYZVf39Xjq1oPv9xnMgLZI
rnwh65HBmd9gY3ECT4TWZ7sN4WJktZzQfpN90Y0CgA3QavHmmpx78Ez7vKItoXtZjvOSL33mEPA1
VkrIBWA67/PVzw2U/TKcYZ5WovqLUCpF/C2NFE4Wj4tLQxLYH1iEoNBPEoBv0Dgt/tCleveEl+PY
9OKW+TzLRzTnROoYWhi7B8nAaUOp2S8iEjQFNRNqV6q9zst2ddyP/LjxHwrCf0iJ21qsh39Z83Pr
vhwrjtMuoxBrrGPp8tbNhHymPEoKu9JUimfvojkQvW93O2y3VBqusYQiLrOGlvdA8S7pQqNNiA8k
dLSF4bOyf59MCuDddnRulELp5npCmvycqA6A97c6K51Jwrhr8P+lnO8LnwZ9AlLzABqzI7qT6kcM
4jWViA7ckrHn9/IiMKB0M+DeHeJTGIAPEakq/Ry81xl1N6X5XkLQSckL/epoKIPPNZAYyhHDxiJ7
gMeuBMm4I8qNJn9iq5qdpQjU/ctgUPqE7sZbKSwjpPcwgG+zxBjQJ3sKWjhMMOKnR15Yk75lpXq9
FDCm0visYkE2vnGMWXJj4zOQccUd+rzIYUD01VgxBWcCEh6GNZxpCDbVxzN0ZfiJYg2hhZKd/S1I
3WLMMcJtqzZeo8+518bABfuNvoLcXqoYI6GmIgckmnk91wA3YXWR20qyMQtTq4Lv5PvMO8Agep/g
zjhid02GGeOeGwJzhFFWA9CmT/ey1T/Jaba3CGWnceVYM+LVEc7yttpdRMJawOYFIlKpqtzqRqp2
NtaOlazZAqXijhwdprlfMds75nSx9JtvBuG49gWFtaJYfzCYwXao8Nuv+EiqYxRapU+FQRiHlcrV
w7qQW7dEDi3cKN1zKJuEZlNHqkaP9e/dDdPtDg6g3PlmsSZ0RX/wbqzqJhU7fsT1qnhVbcUtfMe/
GiC3kFmHgEJv19RkZpgIqgCSoyaNLZ3QIMMOSN5SLF1VOs2Kntgk7Vg8Si/iR1NLCxfwthrAFqKr
U/3oQNhYTF1/rLpdnppolTmu/9seh9UjUGM+540w+k1tEaVvcZggXQ8Q2jZLcpFLvPeDu1yaU7S6
62B7nxTD3pawQ54DKJOsIX38u1is85ZePbQLCxz6usm1VchaWQ5RLg/+snwFh8tdpvoaFT9a5RW1
e0jPLMknBx1hPMKDQbChYZ6519wljMq5PvVEgPYP5OsQeJ2U9YrbHBdsyVqUoQ104kBmNlDTP8gZ
qSGty+gl7RagLqSpzfsFtdzyOST7l/mxJ0PpIhd7CIQ5vzYY4ao9V3Aa/iJyfmgQEUWxsYR5wwOT
w9yws/XrVtdo7CRzivABMV+0KNcwz0xFxA3wVOAdExdDgpAP/i++Dw23VHukMR53WMgvaTIoL5TA
oY8xWsZBP06z8gGQabj6BunjVpKH4HslqeP/jqUglTcAl5qgNxjQ951fsyZJyHjxqMTDuzWBF51x
uSTEgMERmxYPWCoKGWJK7W5p8lZeA4/qrfhmwYdVWWBhw4LttgjoqZG5lJlVdtMaLGQYsULnFSoJ
0ECK3U/LWlGmQlqoxc4KmIa2ZPMmZVdUNGDsRFwXHbHglD8mpxrGno9YzlEdQg+zI3rM7v0CXkhr
PYpUNBiB1Zh2TLGI7fWiWWCgvVdipJGN8KqErVeKfoQFYX+ffH4Wp2KBr0dW2i2vVORDtCM8fdg2
B85+N99MHU2MlH6LzyZw9PfYspPjyZQNzTgT6sly5R62UE0oLtTB28qam/iyutTlQKW8QjbkHKgO
PeKBLXi4R8p7W6gM6GblDITlClxHn9tMhMaRnbkApgKo3oNDEKyT4EoCDegEnwAYPSU44APLTTeE
8TgC7kv1Kwgr1TABP/66sE5EFC9Wb8x0t3T1G65ic3CV93OsQl1IKC1P31re9GZh0Q8qOYYh/CoG
fcENVkLioTxYXDfgh/u8Pak5/oRXBlIzguS0sNZfl+HfVkcad4Hp9FpBbHrqo/cZw/BjF1FyFV42
CKe5MoY/xQ/Fv50fR/offCHj4KqCYDrdxIw1MMYVBfU4FMlqG0ZdmrD6aNpkl1vUlkbeCuy7xmqK
uPTM/6dvVk1tc9/Z03ZSJ8rDXpMe+eq/URxzhdDO+ePOKSIGBiMQKB614zpaCJtdB0/qu+x2hT6r
n36Y028boBixc566XrcUdnV2FrFs57IcZIREDgHti/rGsOYt70d9KUJk5OT/HPQ4VY92T/IDmBKA
JDTbYgx5QUnf8f0F7ohXOjxDCbx92kYpxYqkE4aNNKU2U7AULzqP0iepWKgYGQXuwqXKgnvJ8zQA
5qSnhIE+haURClAbRlrQMs4uXiaN648KKzN50ND9G4jOFqtVLFwL6mkROZD+KJVLw0xgxV+t8nrr
53d0fOUDSbFd3wmi9FVPRLEyR2th0Sbllnr4Sst0P6br2yhTKfONvcVAXqYIMrbjBnbWQs1vG6i1
u2mFcObBwW3hqTehDEFvj95tBgrcOTh9OJMNN2zY9k/AY6w7YDqVf8f3+GZFgNuO455+GXkjekcQ
vJRo4LVCo1RcEDvoPWTZGA+t7UzasDmtOu23qbk7UjGccnhlgnwy0x63SzoVG+VZDn1JtOG/6UJp
pjTbtsCUqbNV9NIFFGim3eMRDFe1i2yY1K4TpmaIOiIchHFocWRKsgwLlrkIULho+K+wYhBHZGzA
OmjSLhw7G7RTY09JVbmdpkQk8s/jvfmkrsYAZaROCF3wD2vuybNEDO1KrZnNyc/9+CKnYdpRjNod
Y7Nl4wBdI+xFcs1Q3abBjjTuKBBQPeJkf+o1F1jo1pdr2ZMvgGnUVRmbJCCHeHDtEeGhI1mYhydy
CO86bEJZDoPx/NlenJko1VIr48zaK9jk8utUfGWD+fqQ3Xv7vo2Uv2a98CR88f/K43MjNn8ywAcR
P0c20YI0fz8bOHXok/sEKBCfl2S11K1v4Rle1JaQn08p1GoXyXju0wh8EmbDmbQsXb+7CRUGxmj2
fnKxTmm5+Tg0xYwqkFJNyjqejXjnJf/40+ESUbjP9DiyTEuqth8R6lGZ5Qe2PQR94WzgWFEIAgk3
eM3jdU/C1PysBMgKlP0HGOSheoZdSx4qqBCEsOATYnPUxItNnguqQ6g5bAfBVSRqkZ/eTKUYZ1CO
H8IpaB7NzSDpfHKGHNr9HTEZGXWZJfQWgGVFf7RKeZ5QI/w0nLyof+ed+kg9U8MVtC9L4MKb9HUM
U0jexdHDYrkq9C9+Z+qPNTxLaojT189Yu7YppESSe5PyXTiT+whjhqruWbVhW3nbdRiiGuCVq2w0
r+3o80yM6rzqsH6wrfyu6cxK6zhNwJEB8q68q404ktkKkto4NVk4LiIdtdAI/o3gx1OzPySbwE5s
+F+8rxJ0bl9ZIf3dqkSKLU6wiaeNOxi0PDvnCTzsRE6uX9yGBd/KgkE0lmiP1e5Gl38WFZuotXYT
r9bZ5RgIcUx0Y+r9oPBiNEzLm8SaRxdw21bxBWls4axmanLF2ctiY+TX6dvRUahQ3QRoc9DFbcpq
z7Fd/fbo0Ow/uB2OZu12eBbfMyMQTQnxynmP7xVaW7lA0KLrzRM8LJHQVXE+Az7AHNBlp4v1c7H8
YtgFZc3dtXVdp5mWLO5BwILJFriheH5VNju6e4+Lk6uK3WS0StZ04VqxgRojqB82p9yKHBOZuVb2
KoSliBzbryi6WfGdW31enSaBbGd3dvzMFNR9/mS46r3HwJyDLsEB9psd2XGO2FpBSsE2Ye79c+cx
uYmJsfNTHUkD2FK3Zk0+qg+5q91WiFE/N9vUTZCZrHAiDQPFZ4V9dhJCBf8m43gahTksN5e55b2p
er1LW7nkGiVZxU8T9UP92nHOGxKsKTKAKZour602gaOEoJT3jVYlQfYJVlbvbVTZigW3h58HAOOv
4QgG0SNNLhLt15DvtfoNpJYCmKPaznoRiAtpjPb9dNXYOGDNH88yIbGwjofLaecMtp5CkQnpDWsm
t4Ki+yx9nsnbmonfv95I/rvhFTrYMa9LnsBvFMNF3BVUL7baLCzwyfCuIfuXCZCGvQQdZ7Fx2ANL
1h4dao6ETkI+PmV5sx98mJgEIL+AXNJeFABFdE0niNIbCyY/tP1MZxzk7kqlkFB2/ZNSsJanijcQ
zY/Sf1at3b9DPR7C3EHcp+8sJRT37MnRTUqWbV3LxIfVoHwDSIfkNb/MWhbwdZprnhUwjAccOlDz
YkRNknOooqsYfM4MlbYEyS7quaZGpLEAbjhBIFOuoVlU/qTgCfSnTs2wKBHYSMP5Wg0kBWgKR7nR
JK4SNagWb8ZR+xYCpA+pj7VkIb+GdbknsukJA9c1qtjeed86KA00mOze3NuE2ynIxAQDoFC567Zc
WEXwwREN0Jhom+7fGb9GF2Xz+nOrxLiO1XTGi8YcscMteAqZR9aLVNnkeQOdHrMzZQjJQ0pNs862
KNWJrKwb+XJIgco81r5Rik+OorVNZFE7adENOwWpfvazPwXCme5+Dp9o72GfXpV6BJ7BjAyIsRpg
QVv8pVBqSl/xhEU7ZShZClAtFR0iVvWLYj6ZziASFBjc5HxLXemJoB6YHW5nY6xJn4xUhs4ELxKy
3yREbBnsDFMrmNPoQQeOJ+gz0Fq1yu84A5v3xmxiHbYbsSVxJUZtLlyEXK1gBFxTk+tCoGgE4zpa
+LbwBNJ2IjX6e5hrtLmHZGRlr2Dk0W9X+AwVuSnASvAdLZTpOXevMziaoYtMVldf45JpI12Aj6cB
08EIwOGcqJM0PvRMZdfVCp4OSd3c6GhoZkfenRULi1YrLbmSoxyhC9QIe0A6ms8h62xIq9MgDktp
/mzlayqhmmHJwTpGJq5LyvnqZPs0VV4ADMUrR3B7fUNy8ZvEsJuJZNSyMmG9kASNLbO+DMaOJ8fm
3JSXZpQqoNlUJTuW4T2tJfpyHZrT5tKhd0KYAdiSpad9W8SLO/932cU89WK9aXaduyQkQNLUnVG6
xiax5T5kiNBhcVJBiu3pxnETwYikM3BZfRDz+UlsAF9amtrlAWfdxF357/dY4BeyLaPVVFFQ6eXg
Lt2KDH3E0aAWdKAA6+0aMAdbjFJ5cEn8b5zT0kBcref8MQxnivyp7jyk8TYnSv1uPqJRbERSArnY
MdwEU2jizM+rlr8KcGhoLvIoW3H50lhbFQJP+yrU3kgv8AMxkZX3tjY24E6Xb5CFi5ISYDFCC3ZG
yNoSxzSzxXzxuiXXoDlm8VVB13bC9NlRhi8yvyHfWfbS2dWUmi8uY+gNaS5a3oIewnIxC0/F3WPH
b5Pm5MiMSVi7LmZI4MeOokVvpkr7FrOLGUB1vB2wQX4S0LTt08uxvoBPmqwTuf0cx7/yGgsliCAu
ebzCOj6LN9EdPQ2Mm5SAbxstSWkcn6QLlvxvZdHhAWxcJOlVJh4WkznxnDjy9HkjE+fW/twzAWC/
9vlXqeyRcycAqq8stc9JUlXNl6K4rPbQKXNKFXGPe8OHkDo0F7bvpkQOvaDH+zGNJ8P/DfW2qZcf
G/Odqds/inDGxMuB5HjQBNrbTnk3QukEdPc3OntJtgqS4dlC4X/ghRfTAVmthBYti1aSKsFkjT02
syS8VguUU1WEzw9UIt0pSjbaO852QiDWEIQc9GmDiLA6QUQOMEHu67cUrvUBP7Rd/SyuMnk9fTdq
cUNNb40tIOiU8EL3AXlNvVIj8F03lLCINv7jLg1f9C7skFw2TRiGBs2BkJhZxjbaY0qPBV28FBGG
3vlxmk0XmQsskaBb2mzVjY5JxuRFMhFKSYrMNHkJGhJOqFoM7L+MP6SB1bQIZjukdC8c4D4s9IO8
/0OfOiVqzxlnN5CyiADeMwBsuTsdZsRJO3Sx6V6CqYYQXGNMJ9Hc68mJQM4SNKkdFQkpiFYBdPdG
r/yPjrRKSGpwB1vPFbY3L7N/qIahzXNstw91AAX6U6QqnTLII1sIcRJwv9lpKni33EOFPQe7AH8X
IXxG1tBQ6hFFLlh5CQfFTR1+Z/eVuUHYJwypizUrlcDsFT0otT6IZCBb/Oyh9scg0X09lWYi/E+1
MeQQJ7YbNCfTMRvSZnnQBE2KGJK1Ja7LLZpNWOkbfNYu2nrZij2aSIC4I/D5WUAE4M7wzw5Fjw5l
dhEM0RelL/0iHQkoHOdNxcgdJPaEX0fLJX3PTySXwCK+QnWFM7ogNYVMyjvWUgqfG2k5hkXDuMcV
b3WPvlX/yhm1+CaYQGeJxfIYzvW+EEx1eCbI9QEtY0j1k0O1+ejqZZBEozi7ZUl6CNhe+WIXhtWP
bkS3r61gSSNAA23HnkFuzewHA8X9JZLVxzhh6ea0Y2GF7MOmdroEQkBFIJMUS/bhoLvIF1iNZPHV
hvKQ72Z4ERs9d5FMnhcCYyfOprJ+eKZAb/PMTyJHzhUaj5WXNVQJ+N9l6jm77Or8Eo4+xlv4R8Cp
7e48tbdqZe0PTQY45tMyrTPfDDm3X/JNMakoIc3XMjRYtfRleRnO9Rcvx/sLr7gwe4XhDp3jHMN/
yTg+M5oy5xRsBJX7YkSv4BE/UjY+FANdMM5mvSTJQcPbBNhvVTmalQ61MzG1LsfuH7fnwejCZ5Fc
uh/sMhCEi4sqBn9vosKpxHRnNkdzU5ZWmJUpxqoyNIr+Vios0+DrDt7Vm7JL1fKDDsvZb0LYcuVK
Oj6C7YiLid9HhLWOaqJU/hheiAZUxiMjx8UFfORJ8f5LrWMEPRXCXah4w8OECgQGgFqwSiCEMaBp
m4x3ht4rCfwc9VPoPtifavnvFXhsC+ojU9KXIlU2TO4MBfd/wBuddfCISm5CpuuTJWe53EnHTfZL
jXFwTRP+MOsO+LdGflTkuboAbd9dKzz1aRP6hdj8t6pQawCobErzLfqXVXLQrX6GvgsdRff/7FHr
eTNc7ltal39Fss2+7eTs2L/VqszlT16wF6P3ybkMrn2YFphVScPGdvRBgKLh1jfMurwnoUvkzhl2
yPaMTGaE6V7AhMVO4/VTgtpfgoZl+kxQo7zWrHvcRk02LXlMnorzc5w+Y81ymGlFFPrkm9Bgy3dh
rGVoCEmpfWxG1tcv7zCP8t/eUx5UgvbxozfG91obskuq3gPZoogv8MiOAJNtOclAr/KOyeqwQCYB
6R0LPfnfSIP1oMB47VImyKNHXdOm2xUXr/aea6WpOXEoeQjtbGvzySs3Frbp+gEaQhDZqaLEIVBn
L1kjRf3Canjw7kOPdxxH10IPnbZP1v1DFsFiYJEAjJL1YZpayJzFQFvVwrgLsb1g2qs01L9QqKLz
wRarnlDkjVb3bK6yFeqko9Yxohuyq7OyrjBP7xf23s1e06bGLKe8FxJn/Qhc0C0R8OQAqT96JsvW
C9MepKZ+JaCr8NBF3BAOj3dlHQPbdJyTlY54AXQHI/XdthaHPLMRkH0bA+ZY3jnK74DBd1ePcdEh
J+JqWjPS21kRBEQESubRfchY440VUW7TRIUkkNc32qeenw1nAVIf5/Gn9Y0t3F6498QnbJZEu4te
Bp2Yj4gczG5mkHcncp5jWMAA+6vVsDuM93YYmgRlInksaJeJ9Nc8L6oM/0+7VO6lRC1gxRTXnKxY
LFyld+qxKSrZKIc6S3dVYIiRNS/uM1liJNgwt1skaC85u0d1nM705B+sbCic+mYLE/6ua/kt+NcF
p2ES1QUytOMLqfiMu9+6Hi3WEYw6HPT9k1DRC750iv2Qzf/xTlRUL8EPZSvV7PJv82VHElr2WLb0
7NrMxBgVLt4MFe3N5W3lLaNGo+LLTJAyoPnrllWitdA9Z2xJpl2r1CYnudtfHbeX4vByl41rZZ+M
PvfJbHxxOgY3758UtsHqWHuWB0MaLbHNYSm92aBW+6/lzLflji+7NilnnyBCVr5Vun6FiFJaC0nV
wSpYd00bD9ggWOMxiGAqbar8LLlBiJIt8n09jhVXBxI6tv3VqnORgPKVGczGjvm80xDpIQB95mQb
rHmX/f/Amg2yv9010xuD03tsNktVr9mjLd5g63OVgT258rSsM1FIBUJqC5y380eCRio3gGhghQ3W
XcoSerDGpaslvU/CIzQ94NogjubUwnKEX750JjsH89gC3YJxXOoqAviY5awhesCm6S6KIfj/qnKx
q2psyN1jQ4I1dexHONr4pMZsCvLVn/rcMeidHeWshbnyCKMjg8vsTL1Bu5Kn7+ZzsW+5EAo243qp
bBUq0BRIufeGYFdgooIS1LMJNDOuJKEksq0vpVrJkLwYWpsl2zzW3zb9KrK0Hsf2GeR7p8jo4qCW
x6TFmxI2lEREzbbdEbV230Nm6In+PcziDcqTxbmqK9VZhXguFvZb1xlitE8jCb+yP+UT+5AxElR7
+R7xUoTwatvlDxjmgTFMYv1LuBooxh61/tm0dLHO8W0euSa0bZxRIDcBFVOfxluN44Ga1X0uoGse
lLDSiWLdu5jpWidLi2CmweByVi0KC5iijMEKodIpyFyFVN+55iP0IuF3OOs+LqCf0A2hEAAJxUMI
+/MoEMOwUYKfDHsE5EHTAvS0NuWEC+4FzjDc7w+B0Wy41ZZSkYvMPxVxJbE19c+iDN/igLr7pjPZ
aOLASJ5DsZ4hkzkf7YeGkv4LsfxLJJLUg5iN3apJwbyeJCIbQDYj78s+or2Squ7/ZiAuvYYn4nTK
eAfEXpYQCj29Gg5zJC0VW7CSG2a82DLvX4aVJdl2X+edsKO4eH+xXQxPQa0ZiRLZwxqdCW9C/MuL
Yk2LaMhqzAjhgo6lFCr7GfU6k8EiecD4iPTPP61Yr7oVo2tS5Iq93VmQxrevpOavLcyRhtt1I7w4
FEtn2r1dD4pYK6+/HoeGIIdWPxAdd63kO8UAYO9h179rRe1n/k8FMqyGrpnwh9MoN6UzI5t15s99
69J5ua8t4mSKtxcpjGfCPHpxZ1qJhpCaunmqsrpLYYoENiViBtdhAhSEZdOS0Q1IxwGLXDrf7ki2
VrHIhyONqN5ZY4IdMOCLzMAGMUpN4/Wb6J2tNGu/TIPNB7DOJyen7x7TpdeKLTu/1CWQS/ud8yuH
A9ilogbXFCILtvhpfCBAO1d2X+odAyuBnHm6uYP8vSmwG/rapk3j1jMOzowM+SVf5D0zEu6Kqh0T
ZvktTgl83czDVE3ty61KRDhwULbII/mAy0h8UhZWx1s6b53n0KGzPXqBe8WroOJ3kNzN2XGR5LRz
pPt00FxLm0WUP/TmYaYKa1INgDQLD5ZTGtN4jKIpBgqw+OytvuKxoeGL4DhcqNmEcW8goKpqBLyK
Re2xXuXzebjs0q3EvU7QpURRer9VRFWLGyZNqI+vRtFv1VfzvKQ4a9mdYWRIoy4sgzRrINqdoZq0
0TXUAli16+TSDZOt32rIK1NrX6D5xF3IDedtUSM7GZnzsnCpkbLQgexMsAMq31DC1ab2e96ma+uR
LDKrg1DE7nFAlOx7JpqeYeiaQJ0xzVnk01y8cQ8qWOGydGgvFVhwqRp9SGTG9D3hxrWT4LlvbjvG
OWeMb37OjgB65Qta44yNk5r9ZZbNBpkbH7MaYkBAHBm1P73qNoQjtHs70jEtDiOcIQOodt0+CG5N
DVDzSl4/0C7BfgJIHRoKJ8PUpM5DS8TfI6PezgAcufTYSroQlbGSnqsDnW0DBapIroNCNsgxCk+A
3J+OWK3rMXR1ds08zrSXPWm3hPgm8YR1gBxPI1S2mP8nUHZWpwDvwZd8rVJUbtZNhxO+H0G5P4Zx
CWbRB/RgycKOM7dQVFf90rl4o8J1ER43FH9Coj3pColpCMr/sMxTD1DQ/hX2sI2rIFrjLk/NGLnI
/NNT8kxCv3KTx1ks+c9ZPJsLYobHRd15o37Xyvrw9Y8+tcTz55idhxF6odn5+NB6Z60m4knTA2ZT
wtj9+imfjsLqVRggAA4vEs++JXJ5MbTcEl82VspJgoiUqWkTiWB3dyQgkjdDWgL1xYP2Qif8nrxS
Iz0t4xNnCQrMMXTOB3aizWfjpxPGwiYyrrbiGqFvJJ4PejLWRXUGGoqz8gYYi/2/fcoEV1fsmEG4
V5Nyl/Y8AY/6eKUklWn8lUzZ34qO5nfUhi9f/aS3XirCYBrvNeDxyLQKq3Uu8rtLlzyBusdXQ2Ae
+4Y4Hito71PdP0EsFv0nx7fi9A7FjvfYWaqgRvvBVW/0uLacpAwdKqG8Z0rKlbdJ+UMgBezEO19Q
9t/BmpnJRIYpTc2A+6eeXb1dqZBsAEdwnqG5Yxq4/oAy53JGxLWU9UHz9gnhrznHVIzMqLQGBR42
It6m92lB6atoSRwj5vNFbkM1q4GxtQiwVk6jhi5UyyHRjKpfint3dtC5UUbcKGdcAHDiOTCX/Cpg
cZW/t3hpAh+/X+Ack31PX2nudxw6Nvc88DIRmjAfUD+7+2fTH7DZMdVCjusNzL/W70KCM6cx9KTo
kDUO1qjneer89QR+Fb30QmRxvt1GmJwV3gvl66MUVSB2YC8Jvl+PqphyWVoxAHBYUJ/EXk47Swor
X4tBfTDFgsV4EhS+bcaOXg5f7gKnx+EIaV7OCABXDlNvO1UtLq4qwsnaP1veMLFcAZVy/4PsAHBs
hUHg20B7JC0HotsCc4gLg7VVRGYd2QI16j2PLwMdJ67c4X0MEy4oGShEs/8N/BxlfW0KLua9t3Lj
+8Ed+aS7K/zMUy21EWkx8QhJsXKRiUNIatRdIOZT2A+8PymLStDlyFQyTl4Vun7YWjqCngx8ZjeP
0e40++ha1TDo9p4NSTlhkl6i1ZrsjGLJnx4xFW+dQmQMKtHR7XZ0X+PpAGT8kFmQCfBGsxTmuCUE
ABQKqsBfbnBtQuPGdfLF/9e9X+JsFu+grIhBZk2WKjc+l3EEoZAboVVnE8b7og6Jm+0he809jTJ/
qGn35PR9fDB46xvbbv0UdJeFIa046MMwl/u6sFimJNEF04xlEP9CP0Rh+yd5M5VLxiyMpiRbX7Jp
jkpShqyjh9NmGlys03y1vvrZ1riCjE6hmxuO2Ys1h1brUy52jDBJrfpezeQrW6akNERAcuep+fcl
Sxejz2GVpJpvdzj/5C7X7iNq0YvadcWeU+vZpHivAQburfNiRcpHLgrsS4a3lA9dy+jnMLjWxulG
vl6rfFLBFv2t4fk//dcxgN0sjYXnRv5udqCDhi7c3HedO0tQt3Yw7bVzE/cWpnF3tKwLC57AGJby
+qECLfzUpi2h3HKsxB3noJY3X6XWOClX695hIBOr42oF0YnYwU3exgMYk594VEDqB/SWT+M4TLM9
11ku71uHm9bbc7C/7AZhBD7serPQD8ja4zeDc7zjhzSCRbjvE6W96GUG9w12KRpZjVQ1OBwzXmsK
4XlRlEOABJHlMTEhqjy5AV+JFeuhFwjecN+vRhkHJFUSS5goeqA+aSDtsYIJ1IW6MhlN6aBCUkMo
BvVyVHCoN70So1b4Jlka8/tSZsNy0zW6QPsgPVlDOBno30SNfD0spzUzRWSjUp91kjJegx7WFdT9
OseoQdYnVlOsToPWCdSh8zvgUyDdu6aYomy44Lj1evi0emDqGoSCAOR9HOKSY20bWmHMZfbGCLpw
SVBdmheg4SyLeLlu+85ang2oEaoVqzfvRHi4yT1Y9MGib3AXV9lGrBrShC1AvUg7VNeyMIG4nWlp
+acZ2vOm5TuTODABlCZ1TQpNQkav29P+7Pgi5/59Iggrz1gOjdX7YVj7xjQjfoklGojdUsMJIca2
l958zKLU46byXWIoiTid+T2C7lvAN9EZYLCi/K4Y9vagAlFdBJx7CajOZmhUIWypP3zf2w39OWFz
L1b/JASropv8ANC5Z27Vyf9QvTyC/ZX4jWf/VaUCC5u90N1RrCcgZNddJsDC4fRPtZs+HBPwnNhq
6LTt7b+j7PoYA5OhBb4TX0VtNQWZ73yaURC8dZSTkjbrCpfxl85N0+us/ZAAsxCZz3nCRx0rCC+E
6Cxcej8g3SDoIK2seQEfT9TJNBMTP1ES3pa5oK3FskHSV+ryeJ6T7X5MZVS3VgWrzoP4sffqa9ov
VoBnHLNavHTyuXf6rzqFAFPPYubRC6abYUiMyOjBd88JlRTHF/UllyTfeT0lK9gwqmHr7f+y3caJ
8dCXK4foZLoEv7Xat2zoAfwcZhTWvUxsIJeFjrb6je6lSAPYPOgHV9225uidhLMdpeFF9F94ugyc
eT3xVW7byMZwgRPihtfcDm8ANHAV2KzHtq0U78dwBCqZzwWb+TIbBbSKaGux4KdUN1+yqDodcmzE
XRWGa6sY0xUOs8vL4OzaHNddaoz/p8YEGwrjR0pVOu+VnuwqwI8JcltTLPYKeJ7KbQ65PBopKrgE
zQWEBqTmY3ietU7Ts3cVotMTg1ocVu0YHlcn736eAHD9UhlfXik+0yKCTZyQRTvbeeIxo0EjPwni
p30cLof09COIbeh5bYdiY8JG4MYJq+N05Zby2Pnw7qH9CF+yv6cfqCBhhMQx0ZdQ7k9BlfKF+2LY
B5nPd5vWmBWJTz/iRNaQGCneEB3ZKjgOJ22FOu0At4zxms7vCfRv+hv1LafeiIwM+INCNcJmV2dr
kzRqz12PXLOorMclwDVYH+XzNbzK9v5IGHlRfMH1ayMnWdQxuRPvONn/gNfE8wI7Uk8XhpheXx74
EnOqkDqC5MZa5iH/kkmogqecuFXdp5IDBEKdGmz3aLgJAMq5SQYm4LDF6XFFHa1LERGOdk3bvK3z
ir+D4V6u3ngUKYXvQ9NLijtXH4WcmUiHOkcagc4NrJFL8naGnbITIBF/arzcQl3K9Jj/01bHlusq
RsMqC3Clfl/ZcOwPsEbUChjncOYhJ9o+ipPMfU4gb+bUeoQnyWm4NgMp7K1ZcinTfatOTA59REtU
Sk/h0y4t9ON2svfe1Aogxy8Ovp2/OoAcWxcP4/uEvWOO1VPcmiR2eUDbo/z2uVqOHtflKaRRKC1j
K6HfFuIX0AnHpMc8fsDAmCGm9udLZGSPX5BMFcbc3KLeyQdDg1uZJGCMDlV5oteDJ0GkAc+z1F/P
EELJVtHwJawhD2QxqtUwd2l37kZu3uhaeE8BVBD1OeiwiKew2RDH2QhvqP+gNegj8cQvawiHSXfr
xEXcd/K29vvk9zjDKsKcArv7JpjJwUsJ8U7CWnkc5Cd55ogNvgZ8dfm4UF/JRt8pewWI7q55bvCk
SgOxhIjRZdY8ku3QeyayCKQg92luQLcOZ8uxd0CeftDZoX4Vbb16eAzpiet8eMx/r7viliuGrdVh
X0k3tE9PIB9CWLKvcPvYasEtVxMa8xAIiCS3MXjVPxYcYXJfsu9tgICwiTnyVaH1nEEP6C5Ewr57
FFYupaTy7927RAOb39a59vbv5qZ5E0JLRbNT2xrfF2+EtdPfipEsMnAfhh0Gmg+tVUuf80kovqrh
7E6npF+k30MnByuuV2pRiNsexeAAxyLvDbfAOLdw+9VOCz2ja+gewTgSiRoj1ZxNWEllTz8YUAuQ
dK6gh5MxGl/muVmEJf+ZT5AcCoGjNLj6OtmrV4fKcBv2JwCEouwNJLB/r8I6cAXo7gDsnkel6fP0
jYRcgF4fOR2ny/spmf2hLAWOeEycbOQZe7TjNETVTbYVisIPOIbY5IHw5hvJFCwX8CRQz64bGrmH
f4bdMYb3nWQ0Wl3b8MYQGOizu3t3NBGy6JtaZ8N8+Z1rOYO5kHIe74Nn6FDbz6OB/EmjTXQ4j0TY
yUgIoeIkIhDe6C1K7IO/tqMNle8iN40WdRuDizaqgxnXykyJDFRKGoW5A5PNckXJfCthu9p/8K8H
umL5Um768TVXOkxucM8UnNvwnulcFnqsfcc6ONSuF7+TQz/G8DcqSu+UQ3DEbjEv4ehq/rvDvDMl
4Sp1AHIUegcPi6rQNvx9kswPcfyI8M2l/LJ37ig60hAM8r7zXcM6KZC2HduL12rxamNp5P67ya2F
OoA4YHFcKY0hBfbF0Jt1cn5KtSbyx+4e6+u0dFSoEOASRKACqtpN+jxp+FsBrOUyRh0fq5VKTcI6
G7rLa+iriRgUQSlKR514HR9+t1qj7spoXuBMxC3IhmKV1DwoW1WQfuHrho0XhwwxWv2WblpaGLYp
sHgA6ZvFJuJx689BBwVOlJKKkdPEzmBd7a96j5jUq3L8n0gd1rPQ5EBEckcnREjHfjsFp99kIXhJ
59WGUG+vIMFtB2E9dGEydmM7OLS5bXXD9Gg2tSeAUpOET4bhFLaccXP1iqvD8sydyU7iaN//Iwch
n3fZ7MVoo3fP8Uriu/wzCCESxlLfUNmzOEIckGtD2qmsmpFbe86p6vzaUS6gm9wvF8k0aub/W0jR
Z8i9h+40fjWW4D5gyK2UXU5z7MVrVOKyySjMhwRukSY20zFbZdnkGKiEwWDdAal88p25iMCkgj8N
etLYuzEVq9MKvM7W1b3SJuibz1MmbOrk4DoZe0O1cCzl8q+CNouzOPDOcDmTabL6TdoFcHMW93SW
1K5wmRFGIhUagXCBuRBS5LEptpGl2QQ4ot6zvUginKvTj026aLMAxd/D5eOGS7VGPsz+n0O/VMRQ
oKoa0OF6bfUMqJUkAmpXkYL/UYG4kqKiXyrhHdz5HTU5zxA+F+j5FVRGLuslPsnZpICt9CQMl/6X
oIvjx0gElBmZrAbm9VgFP4NT7ZxmmLR1GPjfbbGW7OTpgA0RN/+hlZA0wwhMrbVMsyYvPG9jwa/5
r2VT87ffpLtRas15oVS76RuRvvyBF2QXDMoosEwpJtj0i9sEkRZ/7UEo9LRH9eNkdeg11ZUcNvVc
2y+mY2mXTYqV04cDpHvZ9NY9Vo+6ckG13DFKwfdez40HbCFh54Q+l0Dm9dm5OQjXk4LqnuTo3bX6
44SoXH1zOgNXK2geKbDJjcarrTLBTvmXw/dTqLrhM/oivvPRDiu141PlvpKbUoRofLDqLeFBVOzg
Y3x2cb4KtoUQyJm2WhcVrBMOzdOiKBw2bndEsX5plFic3+TYEz07eqcoojRNQpGffgHaSpS0w/eC
Bu7QHtUS7b7rbYTCODonpwoCuh6LIjsfi10huCDsxmNLDpmOfGaBTJC1y+fxPhYiFv3RjqF+FYeM
c2q38euhWPDSlUogAOM4yMbPvp5vocS68SOlDcMx1ij2lHdLTHuNRgBphRxR8TORk4tXj7HAUQCW
esSa3p6LENF8SkhGAxgBABrwGPSrKxLMyiSag2XLLgm1DhrfPs2DGr4T6y/SKhHo25N3EUz2T+3U
mIhJzOQpO8WoHA15pqufLrWWG2dBLZ0E+tgImur/331JQ4FixQ3afIQfVwPj74Mb2wdlFlNMV8eG
+gxSN8n1ytYhpUNM1uC6iIqmEBLuPiED5MVPc5moCq65VnoVeDBq3VwcNKju/f8uIzECxYb4tHPr
siHx6bHWVGP8XdkrBb2ifUeNa1c02V1n2o5B4FZnAXFEYq/eg+XyreATkp66rXY9iLl+OmWeTiPH
CoE175kf/enxbPWDO8WrYCuGGsIBisIYQh9IyYa0GPpBeicrDr24PmWu4K1qKKz9EPvtfaaHvEyQ
V4oksxpTwlAxh8EhA1cCFaqtaj5Xw2NeaMs84KcjaNyiMFDa5h5AzF62PFRFM3DeoHtzLEkE/OlQ
qsHUfc83dXaCjltcWrEEw/jP0C7Ly0euLD6XteLeU2W3Hq4SSovJBTW6cIeUj5JIc+L7C6yUm5i7
F8D/miztQY2c4vZh0PW6d5dHB/EBodHkh0OfXYXy7ZZVa/tG45dTre0eruUHFS4UBppyRLIaP07f
+kBpzeyl2pGmKVpu9Clu+742m10ZZCvGu8wvEf2WQQUkxqR94ODiR0wLyGKYzxH0VvKrIwKcJjPX
WfC+FsVsPMmmib7mIAonngQQyy+w1rs3sWV1oYUjKCFJq7l5gUDS4tYi3mUjXmDYO3T9q7wTzVID
A8P9ICf7g4S5D+EXSvpLz2RsypMqrDf5BlK5q8b/7EdKiE581Lf+pkwMh7gct9yxf7LdWG8LJi2e
gPHS4SAuJ9Q20fjXeI/bz8dveP7Dq2gOYVxQpI7SwC9aybwYTfVt6cE5KjInZaFdK0dH1MCc6PUP
abIy26g791MVevzO3HPV1lLB5ionhTunM5fnBwpamtcyDthSxX6Z9UVqojQg0+YryEp3Rn3Cl+Qt
ZLfWgxzJi+mKuOcelwQXpdeXDABL0ySUOaWXe0So+RMv4wo3Qtte5mTHNihZzpeupSHCmhvffTXw
eRCskb7nCzAjXtDtvbh5FlOk6EZTdo5EHTJoSrPUykmVtp5mkVxBOUHZZWfZrXI4mxqWgAAck/ij
Ob5Tn7I0iM4jV3vEVbFEfMHAMam3dHZQ/fTfEV5RRHR/PQgb3KJae2wyjSI3jFQMazLdacRGmR6d
7LJxGyJ6v5bF4l+TxWSpkb/3K6Q5pogp0PijMg7OjW1oFRsrJyvoaVUuEQspkp0jPqv5Kdb17+or
V1oAuNwK2qDsRI8aVaPvOG4Wea6+PPWs+uscuEr1xzV+e1584dhngoeOzvRnrLWHL9EHItC3x/RV
LaCyRVl1hMwvogEGSkyD4z+P0Fm9MEWqUB3F9Ihx2IMjI0Bib+Y4iztW/r42I5HdUyUsWMq8kmrn
g/YK9Z3q6pKxaDS3MXYs6ayjIMJgi1DlfouE8Ud4xHcoiUplhedrFfzTPKvmsDvGZs7bYJqAIHLq
0v9hekNLrAuZXa9fvn91LiTP+OX/gErMEwz5iJ3DDKOqJ/plzQ4kvfHZ6ETRu36PXVyEp/qWeg1S
7CxsIZCxegIYIvcMoAu0azfu5wuyzP5/zGlvBdm1Lf0Avm9HguL4LgwdvpWYJCEPEhDXsSfGuolO
gi3SVGbVpQ9bwwz55Ub9dj1E/bT/TS5iasob6ZP2kXCAnNfPqwAXTNmZ0zsMCaAqwjR6OyKRdAy6
/BYce2tYjmQkMU59wW05V10JtnZb6KB5nQcA87nq2OSBch5ypQanPSm8bxeDG8PulwUbrOxPq8Ey
7Mn4getzR/spd2y2CMQrdYVwWPsDyZS7BzFF2R12U4g0yP/jVQL3utb6rXTemy/VrEyGtMfXHFnw
sUt2FYem1mT9nSrsWUUVuCQk0XXnkHyth5FkmUu33tOWIjjr7jXI7hHKC5W+EZb+fslmwEoQ33qU
GGBHEadbh4DV5d1tsK33MaMX+NfYvIP6r697r/VNmityDQkwFdZuItD/KZmpSGkW+nsNO8H5pe2/
vavU65uwp14SAh5o319Y73md4O4CeRSGv/J/b5z47KOX3LKmInULlcz1CHRA50IM0TBlwboNmi2x
MuGWbWmkJ1RX7aKPi4NWm6a8GRiBY0yGbnhhvD+xb2ziMk0kAtSeR7UFYdrFHnikioKWNsnZUKwS
Ctdjso/C3ulkIy3Lvzwo8b/ik5p0ap19AW5K7b80PZUzHss3j6MqBZ4VOvDvwkQ0xEQ+hj/y8vOE
Py74uh9XmHkhsuAK1jwYhZ2bWdC6IVtmLwb9qSs7MYiXT6tu25POLryQXWvFJXkB6YVenOjkPg5O
JploPvmPm9HknGFTIaEA0yNz4iWlDUoEA+Mm578kzVpV2CfgvuV/ueNOjFZX019hYzdNF6/BgP9s
EHC/wIhyoLveb/jQ0p884h0ZahnTybbcMDZlgiAdNmQyK573uqht59rEbd9kvAzrVProG5Se2BRa
YO1bCc8npB+VV1sms1e1SN5o55MZCMzNJvXTLhUVLHwawiE572/XXKRV/jfQ0d5l9EHyNNQdMzn8
LIspDQIGra/bnvVDzcZpACzyxKCqfAxfh7E4yf/aKyW4IfDJSnKdzk6AMeXv9Yxh7RPvuqBu4MrA
DVQ+gny9LTD/i1o+nYvG+PzHh1C2rZLGC6oxz7yC9vjD2kL88Xnca28dvc8PzOtomUO/EUQFg5Eq
KqhLFW84jmffklKRhRQWKsDGw8JwFWWodI9+ETqJhQM7ByuJay0u/fKlk6zSNdxhNkah6lCLkO5R
48Y9Vsrm0xlEmxTyJuFGF/aVSIITCtGEE3H3X8ZoaYSuLT0w1y5HFyKojOcs/lmY42DIvSobl+FB
iUvkSdJd9Zwi/PAQdNXsNzw6nqCE0rN2PYcAeJ1fP7LPQ8OooxRyL3DqItcFZppFeNtr2aTHUnaV
r33ArtBaH05NjvTFWR7+LnkoTuvr0MBDdscY0aIyhFyvTjacetSpunld7avci8G9hwOnpMZ50D9N
cCNHAcaOIzo+5Mq1lLAPLalR/5m9FWWGUOnMaqNZA5KLFlFxyL4XsconX/LZRsQKvA91ra0S/HRP
Q2IjSKkagj8uCWejiOuBcayNo6tBc+KQgT2CakoBqcPPge9ykW54ySF1+kTx4yVxxRbxMIRBXKyt
eIoHrMOBQK5WQ8QznAJ7p8tVATfDG4fOqYW5QHrMBVX+qRhN1Qbf2xiBzKzDc8TTiH8RyF8+D1Cp
93pk77Vu/XUVoXJz9+K9M/MRRAyHuWEPTB9FkEWAfRibaloO3Ejxrti5NAkZ5Qq4CORsqrPpgykw
40oWK9h/4DYbDhDR2ek15t+dfq1bEg7a/r77PENiyCec8DJGn8bEbSXzT0Eche/BFqAoQpBD7TXl
hsPZdo8t0F4j7m5ZqcgzQArp9D/qgVs7IxBC6WlxMy9UvAQLxGcIsD6yxp+J7AniOM4hLM6fnEQ0
Y3i1q9ukeeEfJLqkBR54Ehe86lZbs4zFcBVmi0MbtojuLYQadN6x/bbtD57QZUgrQaENU9kWlYgN
k/1RUc/zZNtZ22BBkgfgsRLXJ31EPmwnIdfNR7NgCXCm623Maf862+AjZR14UkxiUHIv+2xzGGKp
2qxw5Itq7MxFkIvvxcbnMmlEGEeDVMFnSp/wlGR/9BxubWmNaaxAT4BfkoVVk8fyxtJazHiBjLTY
/910PCbuVjyXJ5iJXmxgoZ1+zfmz+3jFb4SWtOSIrtdFckc56cU8U+JECbNrus08omMYKa0Vr7QM
XJFoQ/Iz2a6Bh++m849NWJ18a14YECpxJKUXSBaQl9eIaYfSoj96C04wNZ3/bVG2/NkwnejKy8ob
YlHEIq0aSXDMnrQl3PrbFR5tb2qOGdJ3ZLIwoZ2VpSFJ3L90IEgAA2d9/By5FRJsgz5MMX3gzMj1
DoMU+C1ECqozhEtJ98MozwWd6se6XKkRQafalovs5wLMXjwumbuW+XpmkClhCri1m7GVM2oDqeY5
4G33yGl1ZMPnz1Yjgn+GdkGPwbZT1a2xdjydlwUksEpfJUx6MfxWkZqFh2YKP82qZsexmA/YkG6o
UVTChpxZs5ewiomm38B0IdsQDTgC5ydd0QIKvP9K7D/L2Yfx+j/Kfg0EMXQr9IjTRrNDbgqWEtRJ
yBCX2soPIsASY9tfd1bLWATTTZEgS8ex0zine+sO0EkC/R6e3eYl2hxOY3jqL3hzHNA+t9Wwshjc
n565htScQzY3hf7F+yMVFsNi0RKshqFlCHl83X30p3tz8emD4+dCtNpfqwLmobUbzfy9D2qLHc+H
5lT6hJ0AZ78ozTa8BmJPt1sKMxuCKI6xr4l/n1LR5z6Yco7/lz5SLEr26fo78qniqcLnuH+m8IoY
b3iw4MLQH7I2UKRlcKhxbE8vqh7AWHrQzn4L2Eg55vHHqk9y4SMUZCGuiGEYJ+md4xEO3DxHfdm/
Cgosk58xPk8UlSz4pmkXpJiBvvkd26pmODNDmkMk8r3UhoZjaHZMmKo2zesQFq+ej6H8dgbOs88k
+dvpp3sX+zUMB9MGXqfHTOmLa6EbV+k8zkt/Kq4ys/Jvuf0ysGbXXptnCz9qEbRkOFg/N7Pbu1q1
99ajd3YYwCbmq89wz6+1PMfx/NkKuxso4OIbbeltQn3fq+HWpmBK3XrR/jxaraq4k3NDmBHJfwHO
NueFeVRKlRk2Fv4p1UrPaG47TNFcdZWu4Oz6YQaEXXs45Qb3O6jP638AA+Y29z3aUQnp14dcP1cr
/GvPsn2hdcCF0qEwpJJZzWLUkEbxcze6CJwQNNGBe9yNcPeQjs6aIQXP+xeFhHzawtiTpc4Wo/8u
EdRuIgQMQFJhMpt0KttM4+dbM7I2nRRu2LGIrDeM4Aho2TLd0yKWF/48aaLM46AMkX0FWTu2fNib
DLszjAABnQ+KIr12qVJsMrKJH8rrIeJ9yRnHo/IqMTR5aXEv8hEZayZwOXJ6S4O1EkylU02h1ND/
dC8oYRL1GWZpp3TTXUCNoBlqgnshrQ1nOGEtyXD/jYti++Sfy5oQJEZY2wqmbTWd5HJ1Tz865O8S
PpHYHRNXbkKbHzLz6RSfE9/2IOecRvEwWbWav7woCAR6+enKrhJbqxReXwNg25kN3e7I/rBsXFVL
oaEf/ksBcjFqKxvJAxk3c4yNqi++AAavpvqesvjJvLi7aAcfu4a874lUzHOoR4afrH/VRUoD1oQz
/E7zm/GYoqWAqa3xifdjr11npFi1ORaN993eDqq+P6o8YWrTJ/7RysqR3DdNQ/w9eY1GIZDLIDFR
2yTiwfxEHq6NVcGlZkyDJqi+h5rNZYo8tZPV2cjKk3qhxg7Dm8XIvj3Lu50Air5TAHKo7DU1ZEqn
6/ICWicAnasVQ4W5vaBu1c60hrzspU0gQT04p3ezAuB6vOQtz8cltjUckiL82rmKqpdaTlWr0eNX
Tj075zPs5vjnNmGiubmELim6+IngHB8BMpLA353KZm1hYQTjbQtSh1F2f5jULCozo7jXQsFvEjQr
k95eZW/m2HxE6ENgIYx8iKmeVFDR9A6orff8Mj6lkhVRBqRgUgsxcnXoptLtaQiQahVjcScUPgkh
eB/demU7oPQ2En8wWKt1aT4ApU+H70KZYNnKaVswlRR6dz9/rAsxITJaMYmCFgNpuasPHybRBZAB
mhU8tWh9wxH9tY9Ljpnl6d1y1wuKakJX76U+8jMku9H70Ut1LSjad0eP2RWtjDEocTe5YCQSfI+O
R4vAFeHWyQz7A3THcGhWi5h0eXoH2jYLH9VStROkQu23f8lK0Tdf4pK+Ng8yUksBjjgBG/9/1i8n
ny5iGiBlx2aLdIsHu36yrSLmOvqTl76DJoW2FVH4QJAMT4pUtqc0E5F10Govk0lqZfQLDwH6RZcJ
LO8HdwVOPhs1BBKqCNLhPOYKI6uxusd0yFOjXxO8TK3exuBfirQ3M+msPYkxSW+yTCV1far65MUx
HG+e+0GKd/Au9uHeZ/hGEqB9aB6MzrX+etHQMmxSqlJVHuNEONooxxefy9vsHYxU3WcCMosFK4Go
D2rfehvGBv6JTuiTZ1As/LG0Pk7xJjEEYeKnry/k9khpa8/S4HICP6dxEjlN2Pte5QfpamSkWWg7
UDqcEOV24BX6n3Vir4bdNqTCn5yI3imX8J6Bi/qzeTSq8u9aJEtbzK9wrvesgPVhILxyefQnqA6G
hxqPKgOm0hACAP3SpQEkvQfJK/gdHlo4aHM2J3pzRZw3m/sJiZvgxuRtbHRcYPPG6VZylTfPFitM
z6LdK+AFkOlt71KAQxGfKb7u92kzyfzYxYaJiyK3Cb0vEGbKgHJkpEIXfW6T+FSpzKws7WYdhPZB
mz9wY68juYicmQ4GZEbKT1o4ERFSui/5sVAojenZTl5xWL6TuDMhlpIblZMCGB6RELBXRZFmuQQL
O8ZZzfczsmEMjB5fQxAHDEYHlp4KlMw6kFP/M1RrLxPO8NGMdLv32kemLAJNbwJJmvO56kMGNFjj
ElUzz9TkQIkYeotOCD5Z8sVX5jvoaJBsBaw1ZjNtAzHcxcwg+jq+fTxNMHgvRIeWGtRe+6xoR4h+
EK5YR6ewS22oOBiHw+LtN1YZfQqPDIVg/Zi3sdJP8k7MdEFVQUdmY3+N7rC4mcM4T+p1ucRWb+YG
rNjIJvNqh319IQ2f+WdU8AdSsT2RKnP5CfvZ3jYMUIVKDdoM2JEILDa8565hJtpIuWm7n4eJ97vp
CUVcb2/5O4xq3fIXt+giFmBLiFdsjKJDEhyEaKa3Z37V8aUVwcfc7nUSAhZJJeyJ4ThsWLjPKgDD
YcRJglW1INFSzFtdcD8/vllMIS/MUdPtozucUwHpWVNohqsghNuQbUU5E6R06yDuq9cqeuez/NG6
KVuuKCyPWmBIC8cTJJLmN/jYKcpt7u38MWN6HupsJwYuKmB+JpvQMxrX37OMVaB0MundPkr3ag6u
aA+u/tzfewVFFKNSoT27MAnstJVauqS1PbIqKIYON7YszFjDbvNv+iHv1DqjA8AyLqHQWLsHm/UG
IKyQ2eeZGtyDIA26QGJ1S7P9aRnSfX6udB5tufk/d5En1AdHMJNgxud32ztpG1IiPyZVVp/i5uPf
KJK+p7IJgDE78J0fEXvU2QwR7B5qaimmvGnP6xhbAeHIfHgV45wfuobWY9p5wSPDvXchI0PV1Myn
4ljTHTOVJ3TFoo9Zv1qDtVfLGhgNAg/uq//zSb5mc+kWIoKp/VyxEI0sxFu1nl0YcfHfKA381s1f
aDc9mag0o47tBZaiJP9x6SMnpVaLsdvjQ6EA1p8140yYUEL85wcf+buvL0B82CKGV5pLW1t5X75R
UwrnfXwHHg+Qj/48atdbiZILappPbp3//1IcBw6PeiLMQDh69qlm3aWUQX7yAnCDLtIStE1qMaig
HQS5Q7AbahjATOLrhDI14nE/P/H3Yt4yWstXqqM1WBSZSxhOHaT15iVeLAdYIDo+YOi7lhQDBpCk
F/6lgzCwzoAUFyzCr3d8WYdM5HltN3uvXVB6/JMLckGSb7qwI8tmVdXvOWDXU09kAA/5Kq1AGnhL
TkTEnFLDzB0FD8C11EZEDQz2tuDPT5h7Bmc7iwpSTT7HqgL7tVxGn7TCAYSqSl9Mmj1w889MZlSA
kvB6XWdLd9/GKixJht5zKjf+g/02mudD1F1fNo9NdOs+kZiJ+wgn6VzZvcjll4co4okYzHnyZ0nF
PwrI0Pkf2WllpC/LyQDooFHRof3SaEIZ/3YLcN0PLGZFniJCegGJpPHGUxBoE4qFBrRUyHlnEizP
tUc6GW2/8t6gPTmYZDZw8Tk1tcpW+dXCIOkkoTFOlRepvH9wBLdXeM7x5ddQhEQ5umd1LcR1ljST
So7edvrTJJJbzJwIKVDEtMj9ZW+Z45DX5yl8VVw1UfQQnXkd3LhalK0ylhuEkWhbIqy8BG9+0mRK
VhRuMzQoHcX+rZWn3dwaZp8Szj3C21+0aML74e3/x+/mpHOzJOEz6c/ASGvk8fGu3eo9EgUBSrsv
ZbRFcL8yqPvp3K4FmM7Y3uFq0QOwHjTD+vF4UM5ym5G+pRp8ROZxOgLGprccb3G9f+GABo98IsRH
spfgG8gpuQCw0+dj6zSILF8/KmmEhbt1npPwBpIsABVyn00MOjBrt6SKcOl/Bwt743XXoaJxQ2gy
Zu0zurz2znQ+1FfMmZ82F1jvW7N71/b1zO7lNeuE1WLrRCKK/VL604+LBVu/P884ZSekhwOrY0TR
NMf5y0O+jH07rF6IDa+A0ZaZH9KgnTCGLpK4fu9F4Hjf2oDLIAqsDNWdUToRvuI+lkpklSpot76J
9tiLk+9jRS4/hCuMykjJjDUSjpnqRWlxQDqnvfJW8AhrBqE8XVg1pyfNOx7o5aklhdO+y32iiX7v
UYdtggN7W6KjASXSIZcvaDbW9/lynC7LWoxU+TtzGIw3rdNaGZKU8qY7AGfolJjzvxp75QD6+b3H
xcTllhWe+QionzpQUugOAMu1QNBTJFwS22nyecAAL36zVCFAqCMoFvmeUkHbt6DAxyDOmK44okQS
4cVkmOxu8ucC0+OvEdK8cLmyXj50npL+p0Pn/V5v9DEmVn074zKrrbOxfW1SFND3Zx79FM4iNL61
6q/iQp2+R7d0lRgs/gAROQ38Ceb0Jomgfn76KpEqS7k/kbBSkUTNS4uyhC59x2QZOC6Q3vNbbaVq
D6wBuapzsNjecohG6Q5L0HWDqOJ5kRmUxDlYqh/4hLFeEeXLpY52L5adEYrAb3GqSwBewCYSqvf9
pFVq3yRVP5oWuQ+xnXvvH7t95H/luTe52B3jdjnMHfFwwkMlgn9anJF+n32hXWm1EDRFvrmVvbrH
h3AEIjbx/8Li7AJf43gBBvwcTWlJMMERPCXlsLYhdvrglvbEFf+a/SHbmK7AM5bviazMtjfd/Ifh
NI5B66BhFYUjC1b8rJve9S5Yj20xwgTSIEmpCkXBxxDWQveZ22FUnqk38aAaL1d8axcVDI/GpxG+
+xHfyjILhU83htxja/mmyEZyThYulKjifX/EnFIfHWjsKF21HnpI3XziyTQX3u2dkVnJwX91Tc7q
BLYEP+dAszaORCgEcSSMQ+yzEqlW2Hg6v1Rxv9rsLFa16UQb4lESNHOjWE0GIp6IO2AfQsjAkuah
FB6F1tGA8bBDxp2k0oJl+YKs1+syr6fEJnd1l3PDjcjavSJEC25SruIkvR+cKMVaEc73QlFKMQqI
y0ORLRFrbxsvJ8V9XJZzQnh4iXY+Xy2EKNfYmgtx6GjYFKfqzWT6SFs1ANSb776dFsxiOhMLFGYM
Qv8NrmEBMtF6gnBMFPjYoRv6Kh28SCWNtu8tSnHGA01Ix2xhGGvqe4NlFbpv1Yfq4Pi8sYwQFQh0
3PYX36BO16NHaqlywpci/ON3YBcgBBoZ+hnA5DKosxPHqymEgp5dCf9RsPiye4sW76/4RYpB3I+t
UTSBLXoFdZQAg3NjC5E9t9GJaT6Ed6QPKj1b0UpK7XoDdDjDkggJaDMVi1lJHR/L+CgdYvyYq+M7
6mCd9SwPEF3yg7wL3BRlxMCCvsYcP+wMovx4z4FjgV+rfEELsB/+EG3JOlBf9cIJqMH06VJg0IhX
kRtMXAXKd4dKLv3wNAP4xLQRuIJ1B7TwUvYoW5+gS34liy4ziV1GezFrMbLQjoPGsNEWzyW7Fw36
8IfXFNwaGOxTTAfwcr0sgjl/KprA8IYeeSKosDoBSCGskt4fYBj78YSggH1fTw12LCPDXhzRN7qp
dtxvv1rs18chgm09OrY+zWb5roJ0wMFIaRnBiHmJvzw24lLezvk0K91y/ucDU5Quz38NqLcqgRzZ
iPChAhmklk20prRWOuq5zpJP/A6vLd//UBYR1q0oh2N4Ou+r+FqkYtBtGteemMwacCyM9HPF0nqL
UZIAo06Hury+NwUyU4bTDxrIHTzmmS2sI8vhi6INSkJ0tHesKmeUIFzrt5GQl5haor5HWFYcH4Sc
zraHgNia+rsZhR/WmfHF1fpffogSKodHj1hH9MchKLkm4zcbM+lm4ohIJ1fQSO/tAIenqHPTRr6T
s/I615D1BbuHJ8CxLYu5/nyM562opz64bBkaAl0GYSg10kK+g4c63WI4QUFOWkc41JsRv74Axpbz
llAXAsXjcKychS+ZsKV4MK3AJvjmGVYEHtb9znQFdEcBf/YkjeT6pbybEuvOXDUFsqq8XLv68ApM
mbJv/Im8WfmWCAjcNlbFt9ji4GbkR0+cOdhQMtbGsQSUU8o02bcugkE/vFmPbRWlz6FQZxKNmDDV
OO+1ZKrQMHebPuIJVGIJ50ykvxs1NM+YWTSQn5OQEkUGXGWX4RuY/3XWzQfoiFSTTyZ+pEJoUEAB
qCNDoRZEWT1yRakZvCPCJcx1czOY3SIdsXzMfiWM9zh3jIcocEUGp6VnA2nLFX36ZRUvuSkXnB4z
YzFNgcWhHT4+wxINZqSllLwqBjirqkjZerxm0YSc3sjpYUfjsent2aKRUPefNfoDDMNxgSgrxalD
apd9EpgBRjSJbWXXpjdUlWZtfv1J3OozV424o68RatUZp787qkB+U3BpAiXqShfXE5uFaZORWLpT
V/s5QLk1ZGhPNjhAUWWyihjawbYpj3wigMdO7sxod5ESqVtBv03//tQ8b/RhTFtc4KTjBQ115zQX
q3X5BW3ulAgYdsvrYGAomZoI+2b8JgoYOKnNAa9woxT3hzRQD+VOZ5YE/742KMVFy+1xRbDVENDs
x3Or6uZQwMBrNnPeJcUrRyr9GnjuTvfBajwnM1VY9v2aYJRr1mKUPu1CFQyE+0nXB1zMuDJ7CFKZ
bc31cEVBIb0ATkXQKQRfUKlhDnso+tPEgui5ekk4UeAOG355ZaGeXFGnVpfRPkCc4cFdEbwvdTy3
gE7aqu2jIErzjhbxSVf/hZJoAX1Kta+ei5DTeL/gIhSsiJV9yCa+22VIpIHC3uZPkce4purnJDSj
SwYLF2R0SOd1SoriWBYisihFu1DLzL/Pr5dvMKtJTDzc3AIdDhzf+PFVadYSoddR+9XxmJuTaLF5
rVL88rfLq8pQ7NCSZNsuuuzCyF26LeyZ0MfXehtF/4MGxIXMD7O/gzCe4TUFrdJIAtHEDjPJHY5T
7daz70i0tRArXRR+iuVDz0r93vYxdehLbsuMSsRptDU+2fU6NytFa+xxIrRTObcqm7qz+rs6sOOc
Ommyw07eXsMkR6ooljzRoohMQbGuJgQ4tdGGEYgY91fq7Z8ITMM62hIkb5SIUtHKShbd+KjS+ZGu
cUrOScQl+gImyvDkwWizlJG1UZUT/wcLR6X5BynZWqJ3BIicGlo+FbYC9g6ZKl3s2P+MdxoHMFXP
UIUWHNMdlcpSp02RqjppBf3+yf0UM/qZn17g5gc7TqAOJ6AWYt1W8uMCzKp4MVu9RyIiCfUMNZNt
gQepgfofg4RUVrVJDUvJhNY4UMyD3xVjOiUiOkmPE18nyJrW8TkA/QgfcVW8z1fcIHeDYleGDb7g
0i4OkG000+8N1EvMizi0eSI+aDl8h2tjxeWpRP5GvUy1qEzJDpvTfXl56IceDzGW3rgwyVaWJZ5B
054++ZLJm3mogzlYmCsU2rZXz96WS3cazgckMNuHSWFpqGYhm0DLpRoFLwGeNWnIph/g4zEWNpvu
Vz5jLE2TnhDnLDxnMFfW9/pvuNkrNQZzswMXZl9TbEK9YiQ7ZgPbpGVZRn+Bx6E4kMx2W+WgT8b1
+vR/KqsdjyHBktSEY5HgqGU5JPGhYJ5W/aPhUSO0XLuqjVn6O9VEXPqHRsAaR3oHQt2uEjXk8zJ7
mUlixV5dpwcLieSdILQT9ta5sUE1Sfcj+r44HEklWoIglKNbnbDjz/SwAXaM1JJia0rwNQ1M8GF8
O2PXJrzf/Btoeb9ecmeL4LHTIb3bBVkMH3P6oC10QcUcrZl7rrFI7jq3l2+wFFhYVOmosY1c0sQu
Y1fVUVkV51MTwf1gETtHGrTJZ5TyM/s73Md3rqxXZpQR4ZS+ErJEbO4llGRKc2g6QbRk8ppjx3Dg
Jaeb3N4avFoUY+bxAHZCZDTnvVHOzYEazXtXfUhJtHIUPXcdH07wuUEq+quuIb9vi0izxl1+UzHj
BYIfrMHFDAPqIRvHDilE3aKisHJoddUw7XUDbT9CXnG3/FCu/NUMyALmc6JHqElfn2m5xh21vbPO
sNrnX0OzLcR8XjPh6VU57qjrP0o/RGiuI/LkEkCJIo1Hlw8k1BYPH9F/UHn7DuTYsSdNrMkkErXi
nGEkiFU2TVmQNuIMBPnKQdoyCVwNR+rSEZJlfK2EYseuiIEZI6CdnUC1OtZze6+SVgJuvQ1rplyr
X04hpVlMBdX85bItG52ff+6Nsm/xh11ZcrFwthMen20Y17WqCjtxoMz8tVmZXjkft6lOoaHjqNao
j7kN/cQHghR9MsgdczsfkCWWLY+Dy0/EEBXqoNlDzTOgrh3wB7Z0ZCtwhyMUGt56JvbjOiAcuFVS
iREtHz9qmeYSNGLyOXU511FGMgMabm0jkWK+swy58DA3oZZcWscapXEVStnmpqjwqKbAzBY1zE/J
C0YUkWk1FyhfmaxhjTUmPiuqVgN0YbJNAPj8AlXVFjbU0JPYCuT4PW2CQoGOf9+npjA03SOVvkXV
eak4Fq+p6FyXJ9xGjmT0DSb2b+CrhuFBXl9j08w/Rh8Nzo+X41maYw9Et5pisvT4VRg+YUryoK6i
uJusXSBjz/EFMS3KPPWyOhPzeFDlZ2cCh2dn/GFivAumc+j3+GwCHhqWmF2b4gA6+txub/pqEXO3
G9XWdQjlqP6j9Bw+ztSC8eF9/vyd+B4ovUCq6pUsjt2F4omdPLjYRASAzAPBCUqkOvfyQ3jrM+0w
qf0Da19PwKNyRJJoBNKJulfOXBltZ3vhKTGZQWIZSpHX/j/2i/+eAGo+Q357IPRhq5ZEI1W1wo0d
rmbCB44fX4k/W5nRGcYDhmaya0Ncld+2nXyRHNEv34bgLks/CDLPBar5ASyC3n77axmWiOBzRAYA
x/gxPlegu87hEwrZM164vOJSSxhrWtUxqlhWQ/t9O26lSPQlcixvv98PKNA6diKJfI1xqnN1qp/0
6fZoyIekvqGUnfsdKDZ2RM59C62M8PIs2suAXqtO4kDdf6nt3nY8kiRvkA89pHWNlqM56AYkVyAG
lfCU71qqlLW/+Bme84rkKVBqS7abXmBwZH+UtV7Ks7OtH+41p+yUYW22iJPIFeR26TuaLVC+/G3Y
t29iJHiyZLLK1bwdo1uGuu2ee2+XZhm4ZllYgthAnNAzK73J7FVzauV0eAAO40SpHWIidyaUnsWU
WCk4vgyUZyqKVqwxmudVyTZj2i18ml/fxvnBqES4s0nvAnVzs1PLydN3qfV17uvXO0E7Fm/b6fY0
nhuZcHPEJ1Pii0/Z+PVS3UFZz2jHMFOML6N0wIEASYaL1jkyuoLTwMk+QuR73QUMBOLgvDIZPChe
Cp7rhSG8mnxWbfi6oEo0VP92Q3Bfnv3R/IxagaBQTI26ZRMCclJ9mHSQ9NOZMzh3+IVbyofbVqWZ
VTCXrkxOYddBF8H2cvnhx3ZIh6kqIniu2+Gmi622WHJHcZtxp/45rBeY2CJZ5DOhi6q9Ev/iBGOP
EoNTZP4vAyDhLyOv1cF3qUWeg5TVuoQfll9I4c4nayGYus+3MDrt9V9jt/qhoAqywS8YBuJh9ILJ
tLE0cxRjtqEH/E/QQKgjI+mEgvuiOx77QwMNwBMjVjC3HdZn4/UftQLuVvpsYRuFkhohbYLd1QEy
yrMOGvR9V0maW7sD2lrvI4FyM6EomMEFCQ43cZG8oOi0NEQzYCE6cdxBGoUHtM5gaN4CyeujYqLa
DkYdSHnEuzx2n0ne12UHhB1GpqyELn2vwXIpL28XsUf3ZSETPVjz3pqRBlJ3ktjhovbOuh1wUBmk
ie8zDu03qEOGgMlT8EZrX0VMDThgSpNM9O2flfgKpJLPP+YJpjTfPFTNfjH/TRq054lLGYKPlENz
u5ZTMe8GEFCRIDporFWoJhVXEG8tildgeXLW4JvEdtE0T9lg66AyTEUKNhA8iEO6RsSEFE9JTinz
mIp2yXgLYNCBJU4zXnWuAn3pLOe34yJm/gJ3Fcb+JcALktKO7wZFv/26zng3UGOemdABfHD7gYkZ
ARqBCpAAdjlGwSuFSqqxPTgqKYNKZasAGPIo+8o1ZNdSDxGY8Oe6gsoqdV5rHDC8kk72W4/osIba
5qBh8dq9BUpQY1tDGBz+uAVk1JWbWz2x/7s9Fy0g1emhs7gfVo19e5coQVn79lUfpXVDPBWP4DNe
lsEAZ2wk/sH7+U8ArCCNsAYyHjc1H6hnkU7GxCUS78Qhn6Ljnaik3gvqjdG3r4dmIykLswjrypFu
8UaFrAZq577fmIVDE0ZqQEjTu74hPMjNFJo0nzszOgKNYNH/AHvJyGMAI9DhVvp4XAwjFYvZADxT
AmlOSfCB5j+wK8T7QLQC1BEIK0VAA1me8//YWSWB2M1wEqHNL0f6o8pBUGppvIqBDXjgxGoJ7DfN
KNGKmWMYeCeTjTk67YD0VxyYVNQQdJPA29UbyE12jOraN1r70TaLa6E+A+0r3KGAcQVcUPsDbnV6
+gJWdC81eCDo0IzoSu6SOQJW82GV+wFMaGv6eE7v7CePF/C2Vm6jvws+OC3V6B2iLPFy121dQvpx
tK8sVYNe78D9ohFosSscJPgv0lrelgjPqa0kg3S65/7wmz80wSCNf9erod98JCvFe+FapwdemAvY
+fpDjo7bZ7VYK9Mgb3E0+EyX80ac5xInUZd2UgoUyeffYACBEU+00N20ZgZ/X+sRoJf2YjgZTnyK
XAfXgG/BW2fAmboObb7pnRO+EkeHVMp4b1THLdd09aMxoLg5GQqFcUK7cIMuS2vyN9wF4MFpDQ05
QyAFikeB5rexep6X0M1jvbELjvH1Kmj30z7k/KSIeyUb26nmJzM4EeQ74cXIhxsrb/XcpD1wQle5
Q8MlMX7jEGERpUBMsW71F39cweqH8njb7s5r9axQYzFnQGRL96ySEcMsrfQEjLCmVm+yClP9C41A
oCALg+koxfiZ1qCJN2ewY/3tNJEUxLHFa7JCoAoqhPw+eV+eyxoxsGI5oTBsY81dPFQF+xmzC4T2
HHljW7sWg9CBAb9MSfnVasNeRT6QLojY6OoUzGKp9LUOlHPZy0PBuN77wtGCy3+7H+YyfGULGlcf
WazgRko6IVi2gzwDoMHRtICgd7KEHMfbz4a2G6TsI2nC1cOaRaXbLscdOu9Hw0lwjaH5dXjnuS05
fn37GqYH7DTIwjWPaVQk9xEx3H8EIadyUnXpj0cYiiW+44+5GMyLqkZ5gsmJDd4us8jhIeqYYpWE
i5irxbog1fNvv9qsPrtvRdxhtNSV5El9HQ2kjhXoeiLqtBPPnn7X0iq7UyqMEZGlm74yGTKzG+XV
dTnUuD7uKHI97sYG/Eh0QjaOV1b8Nyduds2JoL3Y1wWDAOa/pK8Qb2q2ouAHA/5HW+ycD93Gp5cX
QctNpOlw5ZLQOQHY9KHJGnlpbr/+rr0m/AATHh9MVXWacNe2i3HspJVu3gqShP4d/ZxutlSmkLxm
ufsZ3G9K8yHZIC8SN6ENag4erx1Etcalo8HdzZM6woKsR1USUVMPJhDvHErRuT3RVR0PzBunvD5z
n+axXBPxvR77UhIyJKgrCujKw12qWUkKy4XeBjAxgEn9wJE3r2DG6NHsPn6PULWQ8a8c+2yqV0NC
mzxFgLnK3lsy8x/lmywF/jlv5b6vZQbwlWIdtXAvBQ2yKdCID94bF85nvv4ZS9va/aB2HUuSMs5F
WlDHtkqqNqTVlh5alloz9a1IvrtztiaBiHMep/6hMVbtr7jZnsm2xvcsWUZUS4YUJ3SaHNY5wtp9
y9Q6uJyfRaV/tk6L7ESU4DhGVB+RGo3agJTsaU2UCRFTv+FG6pV1CaFomRtzmrthyTfeSXOMx8uG
lJFOSWp3m2XlGyfsQ/CC13VnyU9IoI8hothbyKoG3xP/4oT3arVGnXLNzotIKLgFzsQTIBDxzvw1
h+AJPV+l3j2hCx0YYRLjPxO8Uxj6UEsZsm2brD1XPaNjwyYFdxptIlXLAeX4WCK3tYYIwZJby1Fw
VYP20wSK+o51rEBbGWKv+0eNDmOi4bssmrJ6h54aAHeNhYSg3D7S6wAC3EH38unIrtk0nIRm9n5t
EO/xnYVaG7kvnd99W3Pm7ZOZ4Fj8IwKyhcb7Qn7KbKlsmu76w7SMmQLE+5NE44t6CWtVGX8Lr1pC
LmgHZYyjKTkEUMevjzfiCbA8Yywb2mXVGxfuKQJM3lOrVgg4OzcPetw/DEOHsWFNtOMdylm/mnWH
iVGrMWzIkT+E286nuic2UXwuvUMdbZDmdXT89iFNb47A+dvc1ixi0CIveXv6OxY6YjpzRoeGrLks
DMTiyXfvD0dv/x2mJVY03hxJXCQNPNTpFq0hdHdDUWSUDtufZ+YRT1RuPtOHNWzsNz+683XG9WOi
zt9i1lQBUJejaXiNOkr1rq0LNsusZYxCYC7fXCcewrrr4DQd+mFF4GkoTUuuutQ7RoQL+IUilO4e
lwpzrdYGY+wy5EDddpC2/tJIiGK7pSEAlNXw5MjAUvEDP3N89bOQ83EZWPMvyRMUfcFAdEqqmXw2
/Xy+6LTGkoAr2pgqTcsL8751upj8TYRpmljCyV3D93jMZTtbRJ0lX6SunKqkxDg6lKOSNS84tsqc
9Puz2WxsYe5/hPZvi0ZssKmXm6GzrAsb1cC8B308pdImgkGCaf/eJMEZqZ4DxP9kKR60dKuf9XKo
I/Zg+FuPtmc2zTf01m0RtDwLssLuzc7U8GSSvID5IQ7u92yDADrtLtRwnjpH7bvjdAOuudOPTadM
v2SIoKo9Y0pVVdk+ACufFPiLisUGZ/Gps1sfHMsBCBE3w/og3SifFIZArUqFtn9eoNLx7OkNvAOE
00YvwVMiLk2OmiTsVlmJyjqbgE37W4grNP8B/jfi4ELjWJYJELDWFWQbwUTwXSBHzpxURqNXBXSF
caq8/QZAqy2mOPKuBjtzjySLorXcfN+jxHqXAuuS7x4gD58zmGHBRNE8U5pezjSTdWeu0dQHpVID
03t5tv/mXKwgIj08+8VmBWLgGRRBXZNiYdULZhFo+QRjWsKFAOJQbHvSX4y9h0UISx0oIwERgsoI
bwSupmjF26ygop/jWaMwDDgKlxtandYlPonNQNpVTbXHliYVjUJEQp6xsSqxGPI2bqwKED4OTe5f
femb9YTYrQZ4jtltpmwe7rCKBKesjfKs1cGhKhFkojq/c2gKpExHHCTNzsEHuFXO4kpIBfrkhJ4d
8nmyj1kD57G2LK7rLDSUbPoDn4/YOoHr1SeAyFYLp0yckrtiVAKjZ+sZsct26ZI0Zs9TKkusR8ri
lKt+I7QIxa4FPanGX1y4niua2VSmS0+feivv4IGsyT5DcxM5/wTNl8vFHgVKqgsc4/Wogp0Wt4WN
V6m6ZT3Z4Lk4St/mJvXOSOcPTjkz9nxb9j/boxrMTIGa+TW8tJKmjm8cJcXXRfOzbyem9+Qhw54G
NnwQpMuO/pYZna2CY94j7E/DjTi99lewveRtjp6z4z4bfErEJtGaOmDq0jBN14bjDw+GXgmRam5D
u4yCMrwdSRxPgf778yBFhQmzXE302zKrwgX/ktu53kP1zBW4zQyGtp0+fF4gs1ooSqaRS1QCBFMD
J7X5HiHPAv1Omz/OS+0IKil8BGrhdU3+NMU3PhKqypDRW3I0GS85nJssn1TnKaXIjhNCJz6Kv0aI
KeLTrdkllwtuF89RgMLn6N5YNmo1hnM1YbQItc/BMXX25HX3B6Phs3hLeu0j9Vu8VmAhBvif6sw6
HqbWvT6znHubpNS9NM84NHrKf3XAk++Cbl4YTkp/AO6wKbbvPlZnk4vg4H43s92NAeEpJJlkftj/
Ei6u0V7Zpvc+yHB2EVvqxPlcSBipWqFvTwbc65cN1Ame759zqEFpvbsv2UGu2lum4QXe1aeP7J74
Dl0vRBkgJIsVG2NaDW1AUiC+BjRa6NQW1gY8mW2VibT7YkWx2l1IC2/dNfJ3OckfPxH5u5UnKZpi
n2I7T7rVGACSwOwwoP/huOnTBFjSwi1TuYpPKL3utThsvevC4r6pZhaSGJBo65rpeSis95yBuZPA
UbQnav4B+VwUy7SwsBwws9QepBA9NU5exNSvbnuWaS6yLRCl7X6t+EyTrUaAnLf+3nwxp1AvjPhO
zZ/ZNykNn/HKlA204xxqYv8VJhtleRsMcoJQKc8AOMwCQwimiZ2tSE17YyzBsxK1y1vF/Fa7Z00p
rNsYTwzeYPflRnBWprsvjD8wFYBjXF/g79KsG6SSA4uUT4qjHM9QoIYWSHa3/vw8byDqdSUdpA0S
xbcdjPwbRTf5OO+j1y5+zrmWlghF0VZjqa4JXcTyag5BjppbOYcPf2lyTbYc1kdGD26ufN1a/82K
D/siNStX8smKN/PEUEbGlAaME+4GyN8ZkZBBrluWKGbJoMiZBxsdoFHogMt7kD3Jed0yU/OmWzIB
THPHX16aDgjPQE50Mw/xSTiPzN5Iowle8uqHwGVYX8xpv0c5oNwRLuVnQnyxCPz8TE1TRRrP/Le5
vDHNN45WlXvLK9CfICuk0HHqJPUnO2n9Xp91hqAJS8J1oDH212cN8fv06GKZ0llgelNiipd75Fxv
WsjiZNVZgt96Kt0CuYpwkB4M49cI5AFOcDfC/FoyfVpLlfbzDyoVje82B1h3gsc/EdPyIU/VSmv3
mPDFS4OuNmoh/1xP1X0f956jwxOehhGnVQrHKY6N1AwiRFEO0bZACyOZYy4wSko9PNy9CtObCH58
/jWavWrqYu5UQ0o2qEwp2D7ORHZcwdTi/140qwsK6xhQbkc9utQcz3eGav8pJ7VC6zmAfXNFkquC
ElEH2JkQb9cu1NVD+sAy0DnLDnLc2YI+8JlSQ+FQCicfgd8qARsAyy3K6qH95UPVNdJT2DykRrEp
f8CcNX3a0ZYY0SqaWBeeIR1pHvueIOhL+Khqm5vC68Fv3tvCTpiBC/iKHMFdcDkMdJcyM2/2U5dr
6tI8ki4XYgNjHbU9Km3HYjO5tI/lEx9fsC+9rnBlJdfQEwC/VypEsr/q0AuKayPnzvzxSUCU/nse
+gnnVP+AXc49k3SUsKrsoUe1KIsg9UOTSq8FHZ3gBaJWAxFmk/NWEQB+I/8t9WidzqtI3lEBeT80
fl06bQeyGeCUZGBSXHI+WtTqbmD/33UFZ5opXb4O77f7BBgC55UTsJQDZSXr5MyiyrektJM2xYDy
Dc8/MvneSk1skTwWQiayyGYxf66Zs2FMwGUSw2BN+zZuskzMsWxZIKFyaC2TY6HvjpaXAMymypTW
+Xal0tX6P178EP57o2XdbmpaAoJ6HjyVqsPK469+Pk9GFzsogeIM+8tZELuCCeJcfxslK6UHbPLM
hC5i6KzAAJC1JFSsoWIWSYJn0gERBCqvclTyRMuzXa5MSP6yDWMG/m8Pl19xT9P1g8Uc574nmWNF
cMBJMvK1HgcQKrzFd9V5fwlVEZF3RJ2XFDvAnAXhYFruTC1ek6fmb2bNOXDRHZmMlP4WBgmq3OIe
DlCsFei3udz8I5FfGjfgq8JLvSKdiIsBIeWOgGhCp57iPjB9AhL912DHwxBLq+Z5AhAxnUQHdoSR
6U5zmCD21D4UNUu04hMT42cLBOPBpHE8Iye568PJ8i3y52l6l+7ERUFMYhLB/ROtGBA4QzxRItU/
OLcxJfAkpbjwLuMp9bQHEOtONXyRhVURGDjW4Ugep646+/3AapAPfF99KbOO/b0ZnGzNMzEjFPEp
bu2jesaJVQhmpwJTDkUsGiH+NZLG6Fr7lkGUiuO1Y5t0nCh9RBqhi0M5jqt9EGZRQnPClEy4u2WX
J5dVRF0ddJWdCbKgJXvnf0ygZi2c01O/lUmab+pNdf3m1per8e3Erz7+tYtqJt3/Ivk+AkFtzpFw
sH6omP8TTnWxwE9NRnGI3rVDvv9fqLHYI0nhh+IYdOpMl0tsiuuas/tfjQo31xl60k8gaNl/D6Wh
KNdQKmJ5ejRiFyYqe8uqjL4DVLubsP9W3Aezcp+kbCqc8CI3llBSTn37tHl4LL+o11sTb8CznBT2
KAbgQ0Sfk8XORfzJPXWD2DCYgi7zFcZvnBA/nniQ237O5x27cwc8cbavjPJr4ezZsPDbejGTdUKm
lsjhowfFyoC09fTdd9+olGZSA3VFosmlKexmVd0p5Kl/BYkUb0PNaa89kgI1JdJaxEcCSwvDbvFQ
qzcu1uFN0WrHBw7YRNdFuYJABablv7d8yrLfmwZ2NcWckatV3PC2/11k7OHeUrZVnM9b/VbadhKs
Wf25ZR2Md6GX9KqkR6fUXDbLM+rqnqQaGu6fLhlyhIftGG7jjwHBkRrlrPHPMKLGgam/J+4WBHcm
YRbiwR/RsEuvoVHUN8a7Jgtu4Ty+j9lkeeAPQytN/nc+ofbEkT2fpXxh3Vi66JrZU9oOPt72zScc
9Dxu0dxBVxsZ9oYNWHFTZFT3or39/IsGsOfUXOpeSJV7nv8buIyk08CE+H0Ji4vPrCBky2rjfZOv
gwCih1OzRK6qL60zT4k6mmMKSyw5Kh4TB4P9cdX5hNuXzcswm+U8oKHzfD7raSNlGgqIz/jWSxCM
O0W3QZ9PiAFkJ5XUYRbdt+KrGUF6dkK+NhFOuYbonEz7QJoQ6eOGXATNhIn29df1JrIGXZofuYXV
trshHOyuzNc5/8BYWJqMx+pG8maVZuy3i4UW6rQVw/8mIiQKfN/npD9qMMtZLvq9L8dVYuUT2nMf
vjEjXl4THgetk2vsUCPnrJGodAVED0DQc0EgaqNhsFA/GDhVhIG1RlHTo9ZxvyH7h42wh7vzaMno
TSFhLldKH26CHZVfAc5/Mnv9bdZRqQVKUxB6kOr2UnkeuZuJs5atF3BDgyJPHDq8rzNW92hpoVKK
cn653ZIAkV0ystWo7guWY/B48+DZoYMhZcyopuAkZCf1+r2W1aTnjx5H0ZnPc7IRnemfh2lIur1C
Xmep5dDdooeMziDZxwwba/NUdswjExp9wkfeFprTGVghefczJHXak/wqOyHaoXv7DHsCwi4N66Lo
HlATuXz2+auufKPAGALHWofvZmO7huRoV0EtqXGwK0WBKEawwwWSGbZJeCanMhtDRvgd6Upp7fqy
I/Y3Td4JCyaQQ1nOpi2sEVjAfXmcIo24ZMqZxFt3NFfKIAcARX0GeDBuuXOT1TqXl/JPhdK/oMFT
LjmiqyhDoUii/cBdEeCCU/gseSixaK7Q6x+1AejyNeea0HEzk5RNUThZft+u5PjdUir7L4Qww4tb
i0qI+0ODPqW3MSj3DYVXm+b0H1XKaLubhvmvtQEJZ82KHfnoJnsWRhFwTNT0Xg4DQGaDzeWrQUCU
XwzETNVBTrS2PUI40fjkQ7fzWuv3Y/C4WOvP54iyzztLQqUYijsxb6uj9oR/ZMw5XZEVm/dz4iyZ
HMXIFSJns4qLnDmU/SAq7MLrQGe0r+9X/k9Y8wq7UnRIArbtMDuFUzG5UHLkSGlHM0duAaC6tpEu
xF3T0HUuXBBKr+LHkJ95wMFnVGtsEIpmsFPkzPrdx4RDCEKsMgqYKR9vlqj1hS+w503EeCRC9A6P
yDMd24FWG9lDA3sHG3vj9bbUROI/+g9N3raNuQLl2TuVe61fA4prtyiGFLfTaarifBi1mSw3EAdY
PBL4ATu4xCMC8fAr56MovoVQTrRJdEEM9akKXgU/n/ybjAJYjGLiIJXRzJDqobALRokt8GCycHQ0
77a2pQvEFlUbg8CrP6ZGAymi9PrEMKVUqwFVYhhsal02ZsicH0C0VqNIUdxNsTWXZUG8mZdb2cEq
/ZeNOQcveCSRc9rZq0cy0p4f6AoZRSY9GhQVqpZm8zIaHUrrPsJQfbAOs4YBludO+kHrrczFhYjX
8MGOAXcLBfFhTNFPAUBcuP0EgkQVKTIoKY8xLiptr4pr9GWQspq4nko50ubXVJX3lsZKt+NPSXX1
DX+7Yl6JIx2oecfIDUxH8D54V8gxsQY+GN7bBCkwYL2J4K4fQuQOZ0kyJfh79DNfRrIBIx7LPx2j
NsKtW8j39ZD3jyvOIfAwloCStwGiAGCCG+VvJBJMe4Gk3gaeg21HIwIrcuOiAmVSNM1h3H++aXOn
vDFYNP2bokZiVS17kxFBsggkjW6SwGGTrTEyZ9Jh1OivWtclBOUHx9n4pD3GVYV4PpIoMmbPmIaS
YK8k+KuY20yTydUKTK8MrKGitkfhkKwut9JcjmZH0IqZYDjGPXblxXSYW24nXiqfPMnj+bEg7jG8
Crmp7iVT0x0rOErUnDFbckDQWvxITzZI3XWoTyXJ3tj6k7pTrwNVSkXpHiuLP3Uacv0W03qNKh8K
6ZuVsM+ZysGizgc9Qtt5pJVBp1uZgJKKoB4T35H4cKfmPOx3RoEI91ouoQzDXsTalcMPURMDXOJv
9OT5izJA8jxn8YFzxC09ZKa3VAkgGSGndonUoW7OZXn2Z7CLeRlb++2nE+EjybLz/+g+sb9k0zxa
fE+6OAg3p5t4FotCbCSzJZoaifxZ57FVAgseoqATw1GAyUItndYYQdbQutLbFyar6GvmvAaYqCoa
jYWb9uH8ltMwftZ6uUQe+ZnuWS9oOYo2hGIq41y/OekzG4QM3u8gwu/EHZVS4oTLF/S4m7TGf16D
XB52S0J8iNz904vZA4v78wVbSC8X1iFzngjvIQowJ202aAI4EpgNuMjX2bSRi5o3VhYhGEJ8s5KP
yKiOhKDmFo42B/Ie4A7cg8DAOcPdWLqrKZVY0rhh6KKjsx6EZMKzCYEBHqdN+TJnNl52EQg8ENNq
Vg60bkHz/17xiMdF3RlMBe30Abw8e5juDA59f5fQ8zZOvS1UDwouekbRGrm37eHbf6vBjJl9Hziy
U13i37ectNzSIkyJQud5s9tHfi1rOqYcZ0vkNpijGHEKRHIO/F9PKEbZBIhiX6yPiFYVQtMtDTsh
WiRw7xDBurDHsoPkV/CLNorBe0JbZYjxPda4eX1oOqpSkIl/6FFEVqtD8hDbgcm0DKDaN8eoeyZ+
kVXF8JEFQUQhG04/P8aVcv6Ao2Fba7wjNVh/fYEbsJv6M1NZbNUXRHMr5ba1Ylr/d4xRhXOkocWV
l1WHxOyHHJkiWcaKw5vC5PK5bJf7w9G1y/sWlMiif/IZevdgZAF+uo0eRZU90WxiuAjQXXN9uTLw
ykWNoXpUOCfloY1NXW6HxVISU3LdKBxjWmvCcIyLTk8RhqE92rBsLoi/2GqqFO8/L2yLI2kDGwDE
fGXmcL0yrHs5yDkqiiJw2Qnq6DUQ93dLPpc1/5NAFoDb5Q8evaWgjg6mQxIHoGcpdbrwLZslvsN1
TslVXP2TKrFIlhauINXu0I04UPI+OhLiMLfdO8EE/UzbCXEoKVtOP2QV0fo2KH15+VyS5HnXFLFk
Kuptx6vam7qtrsrhfwG3+ksa2kAU/IUB5S7r/k4CQDZlF9+bOv1Y6hNZAH6kAaUANDsIjJ5mFDTj
UbaVEB2AlVhrncS9YrzigUjvGk+E9TSaPIjYuw0wEMFh0fN6X87Ex6oxm1Rq2+N3GNJDK6wmqZ/F
eCogfCtUI2YvTzKo2vTIDDCMxjNsCw+1GlC1PoDs4oQsMKncxUAhTSc8nhcNJkrSrfD3aI/K1QWi
2lBoTldXfbFdMS+B8PAiOvigC0KpktPUazbpNvWxB/DxCwbq4WwXbvWO9Vkg5k7btkVZofdHvwl9
sNus5q8zsGgczWbq7Ly5/UfWyYD5Q8eV6f6xXikoyuiBH2PeDQmbOYYM53RULEEG7i2Ou1j0ZiJZ
EmbRr14MNuQdapRTA1chIX5aRcRvnKdMf26KorMsOxOh+R4+FJFFP/BMMUjFiI7DT+fVHva8DCGm
ZEB1Fcai6xXEtZcMT7uxdEnR+QRUvWbsLa8D2SgGBKLsj/m1ICRV0JqosiuJkUHKofEjLZg9mQDl
XQWhb76L/kyjFv2zRL3fzwDj3ZJX9pNH5T3Bs7mng1t0MbquPeRoORWKnBR8PoiMQhMd6odu2KwY
xrFCUhp8ucZZBEVP+RL19JxyxchG01D4qeGDj23fGCJcHEszUP3OjWZwG+iZIcv/OjtXcQoNFu+z
me0SG7Q4vA0pGL0kdGOo6ub/ZJlnigrzWwMDbcunvVbDS/fHtrm2I8LxBI7RvCbdeTp0pUCpSATe
skt69XrsaSYpycY3Z5LGQMn79XTkeTAwGonxG1XFzEHvbqj8G8+qOJ6eri+9soWT6seoOLpTWCmn
yqevzPu6GFrS0I79Kny16ZMohioth03FTnqsH8VkvF91eMAJKdNmybE3wQkTJHFgwrAA2flRrhhB
9knM8eXkG3cZHqjBsU9N+pUxf9HyqaJTerM5WnTW5yEf++EsM303ia3h1/S/rrOv2U9bQ6fNpA3h
VsKcXL9HcQkqNWKjC6SxeQq7BCMw/R1ZVjWL2+ZtXyy3Kp9UozNtbPRtnRmgM/86JJzJtrJMr7Zd
/m9amTpEHnEHhzljhLCotZje9pnxZSA+8SNGsPAtwYbf2sfyuIbGgtIk+vaFJstdbXnVcdgYU1n4
yEtAjSNKLZfHcjCAfqYDET18MaKmoXUNKFBrlBdzqEfRF1HGo/731suNc4EzOGF6/LZBszUXt4jH
hv1AeU5ZbQ8v7mFl3hsSHg45B4KkXYGJR0wqrmTHGl46tThNXHcXebMI6y4+fa6rsgQc3MVjhZTI
l+uQn4NP5wsy0noX0ybVLKP+Nhsm7ltApe//cp6Dlz5fEAsSzbKnZc7D3DzKu7iVk2ToBfyuk4pH
Wo8wD1A5gOanl1g7nkDfiTpvgi36BJrR6fXZesefnWRRgNs9YKOff5OF1Uav5PdzUHwESBoSJp76
OyHlE4KB1LDE70cN0a0iQbC02UhaRsCBuRUZ7uCWi4S56Dkr03HN/SjAr05PQUltX7xiUByDCf15
RY8toJLePpnyOIH/Te3uRnJp78Y7m1DMkXlYWKNXyMYFhE/9jBanKRVcILr5F5dgAPIYZvyNB6Uq
2xe9DfCSkkPxh8bVMkni2agwIvYVoKdb6onCFmL3ap1DxwiqaA/8DHMQDIDZwZYrN10eGudUqw6f
pzUPNWjhfqs3BGckYMDOT9jb5NA9YdCi4qypXJpHVPh5tTf0tNrJIGFrJbbXz3MIWTBnKD60JSyR
9vpcIrkhxiZg9cJ/ftIbIRcbtK1PSVwzFOlOR+LJqop3xkCfMEmh+k6R0PsuerkzoKUdCfBRfcP2
5THIgFi8FBlwTdWk+hzRVur/46AxZQwSabAAkpBTWnF0UoTecP7pN+IgUBlqeV1GrF/vKKLOF9wT
2xQnEaDb+5blB9SEQoYgJ/GzhRRLsCKTu0AfgBC/UQ9dxNA32ImmLf1r3azdfz8gF+2ado8fkYHh
MLbvnHSF3a67/PJjMFwHIhTPqdVX8qkL8mzYoPvZ/14I9FQQo6zSlACmt6f1DHUWT1uREwschrRk
bbYPLB+WqaRaQSFKvoY/j7AS4k2sqE+MDze1KzQaEIrjdmeXEGPyAxVN+EmKIYRhzKVxFVRABn6s
/FwmVgXm/JbkUEg8TauHxeYgz35jXdcn2i/g8jE3SaxaI9iZLsoXaxuptWyJbcC+dcJLzqWmIHHg
48lEZeLJnaP+nLAriLxKbqW4OEJxizDeZMx+tMBjhSJrspDqbFt24ypxWSTlVIi8Wl2Z03zEoTsw
avKbd2TWJuwqduNGUzIGPMga7dutLXj882t1ihLdLif8mulBw8bqRUSPzoA0qggxFYoa0Td1Yrg8
1OB4ubLHabBaI21aWDgrq+6a4P2h37e8Xz7uTQa0jQVeU1HkF4vE6cvBJoTwcLUgnDcRvTII6Svb
AHqAgp4gblcwPJQQT6lYGeF7HQFwUOZB9R8lv7A372OXuzTLicu/eiMZUhlTxs5x45ggtVTvBVlk
MwZFFRTaFYgepi+kMG7BZwHXDOgWfrMhMVVjgk7EsL6K4yWVsJnXZVBS3s+pe9np6XKDSy4LOkDw
L6TO7ZmG0zDtjNTs9xXvsKEzwlb4aogtoEb/uSx2CgHOxbr38HAL5hRUerEhYbbixHzoKjTgkDES
/wM7tGN2budeb6AMLufO1ga0YHA8bSao99Aji/slBBsA/LZTSICR0rlE2nZ1JuIZaM6Rgl9fmaBe
QBso2NXPsdBz4N6/QsFn5Bc10OofsCCL+BxwHY/rDk+s8CkrJrVfO7Mw0KXCP1fVCnH58S4arQyt
hhrC/pQ5Tex1DXPvzWltGxoS/wgvVyoFsJjZEaNmVGif1NfN252rb95eC1C/j0S+oD2CAS48OpUI
D4KigMY+hHQQUST8omXX3RIPpsUR3BwQjHwm79OON8c7UCI18VAlN/ufHWWgcIQsvjzhjYvHOYkf
VvJFu+P6wCGVJFbgLs4F67oSk6p0ljTKN84gEv6wcHRwvEQ/Nb535EffxfZaepiC4I+MFhStn8Ex
WAisM8UdeK1sxHlSEXyI2CEtm6Mra7h3S9b3wQ6nNriCWUd1zrtmWr0lOTBr3mGl2tLRzjHq2F0c
6++c6tmYFVyU8nwk0q2y9jlvRtxO4g2hAtydACZ5UrHwteaCvH6Nw1DJdq5WSG/smSb2a1FzXj8D
58gvB7pvftcJ5Epoc9SpaVZm6iRbJeMeiZ57NBs9fXJMPc7OHXCQQDkt7vjZ8GxYGsjeIr9EowMD
DsqRGPrr2pJs9lNNlY71okf2Hz75oUzCB9Ydq/f7z/glZJK9LHRUqVm+Q3NhJRfMigTZG0cwm3r5
4kHHh/KvF6JzlMsuh3avJ25RUNyBn2F1v5fRqu6bxZOACRblNJW9ULcHj0pYwxqjTQz6lkURu+D1
kzOZE1GwtcxICp/X70xvlhDmYJs0XgM4pm/QMtV5tPPG/CBP7cKw71QCggPkkjRiLn7OkSIlCdlK
KYQ+a9vbsspkCp0Gu9rKmoz5mf+zOu0TYi+UAhs/Cb0nYhovu85hw43HIa6Lsxroc8d6+Mfb67qH
dUNAjHZCgn7lgbRTlfoybKHGAXj8owmH3EH26DygBVzR63BF/gMXZuaZ3WB2IxQDsJ5nP4gUX8Fw
Thh6QPBBqjryozVMFv7SsXl7iXtA3eNgDq77OzvhDbJw/6YnHgKiZBKL0FQRiTunATXLAXRlsj1j
oYjvz4plPlGPE1Cqh6XrtUIcYcZApOLU9QsvGeSHTzXa2H5eUZRTeL/Y3hUbr610MyydUtGxjy9Q
U/XkpvheNcJfQJqso8OOiZz74KIWgvBSSwJDS4xWnkTOGdynL0Z3ywiZGrgOjh0Zs9AROxbyb+rD
R5L0UkyT+LGd3QuroEf3PEOlzcndtUEPlLBW+qIMd6/paD/u0FvxngtnD4DqwclBnv5wF3/AtTu5
3ojxz9+5Ngo1CkScuveWEafFNP7Xt/taA0Hou0MRRX7gwlNfeBdSo45JiH+dU4uKpGMAjv5Z9rni
TMgXf0A+XfnHl/NW1G3JZYBk6kLgCmNkxeMTBTUOivdxkCqQG+E1EPB3gzRzUPoCntjxHQ5H/Otw
cSEYSTScC4edZP5mgfsdVnuY5SQEpiIBonL0doXJEMZSEWjHf3DvWdPJ4ZAoHirBWOJOtMKeLGiL
v5UmgF0QpZmV2sT/XKiNwkfIjZYJ7wvdtx3e7nL8+rtwIxD0Ox1JZ6sTBVFYl/UUohYfLBcPeTbR
gB3XSYzsL6dTGqfmRsrTnKT/mGkwLI4bO84iHDR0ZKgvxZHIb5aJMhPA2RmpoRDfmiXdSWCP2Lcb
dVjG7sKWBtp6V8g0zYtjcLDv5/js8Ra2H5HzMu7nA6VeiOmXoXkDAEP4XvJlQhI5k+GMMBCCx3Dj
oogzhM6WBM+fGAzcSkAEn9G+5xt5x7wACPvYjS3miU13qH1ToTWqjDpi9QEfTw150LH6lJd6qXm7
JzSDxxeGQ9PpB1iYOgJ1lnmTSiFourZC6CpAO9fQ0sjk1N2k5uAHwL9QCwfEqmjHVYTO2Zp2GPjm
QOlRr++f+agQKUX3H/vi0vldjQe+giuBgKWHnR2WeTIekl569wbokSS4ukHyb3dC2EuQ6+xnEeD+
XkXplGBG78KTmt1T7SALUJTS67pF0UfRI+4xJ2njYsP1Rc4piZxLFnt2af4NyGYv58Q3SoUtLuf7
Bc7+VY44tQljRIn1nJaIsSOzci9tXWT02U5EGwvbYfS4W2dWzH8Iemr/xsi18NorvfexFvkkqk2J
fiTPmVBiyswyFW6iO58/YAn7FHC1XrfQZbwu4EPHm/Aat3afDkgFpsSYMlxUHz3yMepRVoAsenwV
qHnuzf8HJpw4hWMCov8YYMSONWwdbSu65z0lhayH794C/mpiL32ZYdUrYJOgRh7FoLiIZ2LA7ucG
hqRtF2zSLnrArGt4qtLRZZzfAORnAHs67CPTKbFW3n/NQGw1MJGRgXNTfhzqrC6S5AJ4IgrOzbX+
f/bvEwZO1tUhIY7ApKEk7RHoaIzzr48aEL2yNs1qr+SXkuTiGipFsLi6uZPNOgSFBn6N81PlAW/p
6ZKIKNm5nCUDIw8toPygFyUyjLFKmAjNpsCbXItVsb+APVJZd/IYI8GWWVRXZsmXO5QDXl4cQpTo
32mbW37XisRVHY8UDUoMq/aZbzJFBfxs77Gnys+5UwcBxsFFnunnGjZ04/rSbfTiKOFAZx085Fz9
C/ZQnzFuCeQTBkhaGzDNQKgPeVowomPCsqo2V6MEl6ekQFg60fOod8QWlRA7gTThLxjSeXOvsTzg
B896W61kFm4c5bt2LTotbCbioz5F4BHdR1VGGtkXJTpnJdu3xmw6dZyCGoNSJovl+RYc12pe40NI
bbnohYHVcOeKyKWm4JF2amj+MF/ClmTAMpyswlsYJtFEWIwYIhmMadp/taE4RjlrwG4hYDSFewDb
acFlbGzXmnnvcA9nXAcSZ8yuWWTIzJEeGC+m3L36bg4Nwq1qMt4tNvXMiVT6QQkG+HRBfyiRVFNC
4enoZBu/Km/UeZ9/tQj5foRVKd9eg4rrpvLVefBWLTuLnMnn2AS9NHRfV8Yb2SpKbhBfEsi6Qnj0
aAuIKKTN8pxguXHSMYvX8UOpjEaLHjNrXcCof9bFIEQ27nwglzWdrYOTAuXKiJzmxXz8QoWF+fG3
eyDoYLaTch6sgiRpg4HKvFlEjJK1uvoDty/RDITfqCSphLHTMxirDtPDtZVQlMUqaBWVYuCKo4UR
33P5fHHmWK/bX/kx24l7dNi02iR9ZzgzXX32k+9rkR8vJN6o4QDzlXIv2fmm+dPG3DU4k/uLpyGI
BUAdAdah+usch0eB1bAi/NvjvY/d07iHKW/OwE5e24rBC9Sl6iEoVy2iTi8Gr5tLQBusbIDXPVQ/
kpjWA5nQPlFLvtxBYRVQL88eUKGcs8laYDNV/8Rt0WuYQwGa/AYwIvPi58dUjeS4Bg4YCiq6/18C
C7okrSKZEsB6VDH4Y91swv2YY/Y6QVzYfxPfxUvmbJAcxcxEeSkBdQ/tyekGUfofLCnBtY94qZse
ExQOmFBb/Z+q2Rz53vysW0dOx3ytiElnQUXdFNuAkYdkggUyj7GfzN6mEIX9fTKOps1OdteogTo3
s9eRWObJZlqd5aeu9QS73PFf9MCVtFl5xtBMMuTx8+QXXVd397TgPyAsdhp5eq6Z2JB7BIXViZv4
U2Zj0lnP3naZ+HPrl/e1UzvoPdnx8rMqhJqPIGJpHWh6kR7AmEM5vWCdWApHNFS+ZBr5ODTkmMxo
1jDoWQ25NOZx/WjLnAmqTKTRlkaVG+IsUThQtcvUu8Vwiy75E5ah//Ggx9EQcGrrQSCsjEsjMbhv
GKiBrXhJy3X8G/rKcc+0NPZLSsB2UhCy8724t1oBjFQMlK5FfzeRBsdpa3gqBzh+PNKfPu4G3jQ+
rXzXf9xaEziqA3nVqDwlyjJimX39px7gecOqdEaSBrhRAYn1gkZLRgfoxQz1NdR7PwHINI7JQvLw
qu/XkKq4/7jOA3m6rpOqvW4eixzuMEhk0BvZeAfxsfiLRwYtQxoqC5aPAZyjey4Pz1c/HP797jan
QCDKNWKsEa7OvJQjS/kMabQjbxiZrD98LeDnkF30C4c5ODLaD9P/Jrtw9DMb5dEM8mdhArWrngQW
wxL9JZh520euBKW+GJJs88l6hV+x5GRPglNHMj1lDFQTxRJ41qqtS4owS/0KB6J7CqJvMhq+6ZGN
s4FAqi3uyTlsJAf2JcO9eu3VXGCAyrIA+MBANChpTzdMkjjG4fFyVl/r0ZZvGa1fOqiNtLD/xMLc
JcB4/LJ+opQJWLL+eUxbxf9PQ8mVE7aAwiVBvTqEIliWiZ7tYwQhOA0kJPl/6bKj3j0/STHGARTi
q1IeH4jXf79n+agdEzFfsqrYBH4xG3XwDWiHHEE0SryNoEYxkfLyehL/J14DpO6+JPkEV5l5Vpst
tsk4Pq1UhzBEFavUzSfh7c/dfL48DyjA73tqeGAMIfzwXFpQY4rJFVZ9gLDNpB2dQaCTuarV8lc7
ZPu7Sl4KAg5153jVeRH/4i+zZ5IbpQcibrfOGyCo/GXq/3mmJXe+/irjSjPcNry/Ra2In6TgBOX2
6BhUgMeaxFWfNQneHS4teKz1DlL4BOSnOm8LKvqEb7+aP5NJYR12xm6SeHL/DE+nS1ZymxEWnLnh
I9wWB8F6Qsb1lT/ZIDDgmcLEZv+ExmbqG8Sjf9N4OmqgVxomKLki0eMKlUEaluUpC0EdEB7uCXVW
pRMNdCZXMwU4XSF3SVr2tLjldFXUfwQOGdlXb27+OhSricZqQTQdUktL0iYPzjcxcuf9wSTb3Lt5
pCA6hL+E8diMN0BEHAJy+AenQf8FxpF2CaMMwOSO0Nc4AOCVTXGGyVXH2moXFxHeZolx/ID1XBgI
2bh5PMXvtyHJ41ifV7fS36LPIqszPAnFeKBdjVr4nUvKs2RqhCWHJrgvH0ucdaS1yQ4VGDNOZYUl
qMzq7xccKkoTe8kc7Wwr/rWYmp2ozW3ke668qMpKR9XelLjHHPN5qdLWtWFnwcgUSkIXSRBfA9GL
ib6MvTKeZOOV5UKfvG+ag+wHZkzSysnuSTUXUDmERtIl3xjLLLxoKyUDErs9V6HnPBC10UoDvUHW
38sMrPKrJTXO59ytb8o9Iw6x/nPe81h/rjXMBe3iAUaPf+uVnSiTi7R0BHKeD5n0b9W+QsNQKabQ
LmMZ18xCtMn+SfOiRQRiGnvGi6TdzytelppMZ/msRjRcQjMy5osXbVi+Ff0gPNNNNi+U/XSQqmSg
lXapSRED3hSsvbzejW2cWYXI2Sf+2DtCHN13DlDV/Sa8xRjlZKcI++xc7k7GtCeIpf4SH8K/XsY7
o7iF3ENWszsIz3o5m/4rctdWIwhSexKAL4dVykjb7KnatXsnpT9ZhfBv4U3MzNTOOiIG+LxYZ21u
VRgyhSjwt3RJ3KsMBI87TQo3HNglfZE7XxQr9/8NNRZkR3o7v+a0V8IBNpxS+4QMR2sSaiznjlCP
FLCh6+XLfJDQr5UDRMmPZRCo/KXzIQZigvcMgq098hDujVMh+c1UMEdEWi3BUkrAPUmX6YKD8Kus
uB4GZyF9dZJFHR3WHE8nuTMqoP+db41wmTt40ORb9em6385NkgX1FejOQ3KsQAgSkGax+9DcfOGQ
Cj2dTYqOAB8jQCRZy8/2UZFjWdTucWRBff2JRDC8zOpVAWmdANKQSlw+aS6/k8+I70Oe/wvlO3o/
Jiev5bki82QzdNDz+HRS4nAgXsoWJ7dKH76Lrw9VFRK+edYyyz2veoAb20+pzj1oDQy/hghql+RG
kJQAsZpdx/G0Z+lgedjNjGTs9jYuDs5BRh/Cofu7b/aLOl8v1qt6X8YO+c57H2c8xgLUDA6/hrzV
lwC9/d8rKM8UXBhvn//R1MaXdAEYx/f1JAWCVLXhKKqwmLpGqe/MC35oggK3oo7LzGuKlqzZPUc8
+La5E3sV6AFmeRkDwNC+ZsqxosFmP5hzRySarUTah5t4Qci06Z5ZcdvBiqSWdeDVXZ9jdiNq3BRY
8OJ2zRI0VG0ydla2wmZeKKJ0f0CIEJWAf1qzntlbfjE6hUvNb52kTU+T4gfSt3dIoTHIc41Az6ww
OAzhybXT9ApqjPl2zVHSb+hYmTjtpTUZKIiXhLOC3B39gnrQWkfggxc1rKhsX2oPz3TmYcjizRCD
PSaDOQg3V7BHo37tvgWv45CuZCwwUa9uJUQxMBofp1QOy9A+GtIFKUiiEtNLO3RGruScU2iijk+l
Llj+1chh50yHuaJRDTJSlgaIjiF57zyvA+Y2SENLlN4EA3vYTSYKBX9knFnx54hp02JfzOha+nd5
m8MWE7+mDudR9Y5cxnh1j5jIYnzWRYpLNgIpW92fU12UJH/2mp6Bc5syoSyTwIBAq5VAGB2xnZ42
WUfzyFD6aMaEbHjYj/B/T8Tg/pUs1jyyR1/qLPEazA32MORkhFcwhcRDhihAUtv+/pW+fZQdvuMG
97u9P3vngXhY7F4Jm5UykLIrPLaziF5RasiclUXC49gNEl3fuFSo6nw0haxjJ/bavDbDJc+Kf9w4
I3sbJ7HVAE34bc0shtOQJKg+3t0Jjj9dVJhD6AyEsQV+3TMSs/u36C83L4qZ6hSApURMx7p/imXj
sep+CuntQWGMLk+hwMOwe1L3h7A8RDUmIJ5w1kRdbjb56ZyFJ0h5VBlFJcbchPcpYTkHj9Sdfza+
7vCdjIsJAy19s2LtjHbw7aFu14S8Z9x2xtAYBJciGtmIv7bepX2C/IWZedZGanipIMkFzi4NRHCr
OYhM0lSn4jgz0jsOpOxlSR4TDmJjDySTF2vG2gYCE9Jzbsn93XIizdD1xCEG//0Y063Eke6MAuit
StOWYP8nP5UKJ7xYOCGmVmr8aJlZbZ5LA+tbCiPsyTsWmplWTNBJ6yiZMT5a8eQOXA4YqwdsgHvb
Jhvyu0t1XAygvw4ONv/fB8aFN586NOc7sXENsvTW4AC8ioZnYx1+UwPO5m7eLcYifoNbPyTab2M7
W8UnNTygvxmnCpiXCCo1j8RyhgIBjegnTcbwc30yecqnjykhh2T4Iy3G/yu1CRYm1vxVi23qOrA+
v++9JRuj3nzKh7HsSew1DjDuUPDfWjFP2LOE87NtceUsGeZ6olnhpEih/fGx62ILo6KsLplMAkhy
vfG7mM5scArLZ5Riq/OnmfrJz3TdC7xXmfqX/00pyfvOxCGKLSWFHdXNQiaFMPmoWHq8M+47hm13
GAwomvJyLevJZaTXtsfKXDwvdJlHFgBfCRIm05CAMaraUsn0lVvXlypj1L0HDzvSE3KzbIj8QHHV
LtbtTwVVTv51qj0SijBU0PRHUXohQ0rkbGGDVtXaZTbYBb5c5Im5vnoaxF3RKS5OkLuev4YVGlu8
U7R0Hbak5syYoPIjVlu4Lv6wGBWqe+W7OIdL1sA205/hcX4Bp0I4PJmEFOQDh7k+8r8Oq5EV5dn1
b7RZM+637RCuCRI+xBA3H+fGR6Gx2nA5TRNCKO5acUJtbx0jXa7t0w5SzVdHd4GNHrCIAomeHZow
Vt91WIKajVbSnndf1Qpyg0NqbUpsw1FWL/mpzzhNlI+jI0KJqv2/EX9kX6TVdDvVcG31UvO6aMIp
JBPFpGp7LIbXycx9kvMq3VV2Fozkh1oTeL0z1UmNKgNBW0wJX2y+rk+LCuzhmniNfDViuXmnUXr0
8vNsEm2yfEs0wT0jrB2fQP1LKLz93k35F9G8BfF3oYSd9w4GFMAhxWqQoZLh17K9UCIpe+QUfawO
ScmAYYGNfGxn9WYq2q1T3vlV/WyTW7FIP3qH9MGq6K4JXXaMvSUWuKniE7w5Qv1/LsqMP9HEZdu0
9nBckGuUcHepKkiNpp10FlecfCEE4j8It38XdbzVSueTEmSTFCRkbWVExWla8NAmTJVR9/vXzUlH
TI+YzpX62Z9+x5gRRhhJrNx68P445wqast1GoZek0RwjputV5wIOXxyH5z+PKb0ZX0ZM8GMPiprS
eAS/FZeKX22qDrXh8rU5iNwmCu5Te/hvIo/BmjNZCaoppanW7N7qtpu2kp52R6+/z/jLxj2l27sQ
ASyu4xoy19x1HYlS0GEUYV9gZ9+NEk6fV1K8pfg3fyyr7U5jJ+eqMHPzQnZM+QjU5wChvvcftAnw
hLjW27FerzhUlg/+wdfMjnBEOVKUHXsbzjc/LB5RQzUXAUo79A3VEQ9y79SayGhOi7dF6gonJIOO
usNctInzeI14ba7D7Fe+sBAQI4qy4WLtiABWnDcP4F56CaTFY49ggb3OKCdAd6r4td0H/zbJNoTu
j9LUs15bB472ikZXeEyEVWqONpkmXxa3pOm96VJEay1SdTcBMtq4lPjhGjR1xq+diilR/LexKYng
LbAR28KhMuwYrs/Lale76q3STc4wTFUS/ktzfAGg2Qu6kipSQSTygT08znQs7ooUucfYOlR+1X/C
2DjFTQ1UtyGjQdxlFdDr4YEJDl4BSBOQoLdGTX2plSIEN8XgYQLvnNU4VzsapE8tKTaLasG5xVO6
Z1l98rx/xmfbCncmx7DXEkRmhz8Bz7ncfnDCAzByRhHlGZ+7oqzGpakJrL4p9u+B6fbLjsGC/kyU
ZckOw0HkJhCc6Xzb4/k4yk7h4L2Ck4d4aH7ysRVU4zN5QO5gPEqeq8j+4H4MbHjIFEj850s9XdaO
DR6Zz3GF9euS2oOkWkSwMP31mTdW2Ab5irytklariXEwgScQoPOSE4Qq9u91jwXJNq4CZek/4rv+
nkYL5VI/6jiOgO7/DRLrgbu6brHPb2PoTqDTLLu+lMU9FfrgrvZamLE2bAnIrJhQe1/cNOQV5b/C
R+jyCPGDmAVbFfr1ak95pJmDpifgEnFm52tDKHuZiyJczxtEQ+QuqJLOxxvV7E3ZL3weCr5SHdP1
dQFSjB4slpOT4/244m2hLuRxlZqrCdo7/Gy0QE1bA0ETESdhua67UodDXoqeYq5TndpIOqNt3Ig7
X/qjp4UWDtsdkHZF99ntbunVy9+RyxUedX4TlUTw3+x/WyVKDzozhqySQD99fmWkWBt+xhCCCt8g
5ZlqScK30q0XLc6KTxlZIixT/cID0hqDcYPk1+nC24fHx/b7ufKiMYJSC1h2egWRoxH6HhhvL9aP
X4LkI7v/3SQl/cHY10uNjABKcCQG9EKMbd7wZoFDOf3olE21nQWWvrVHSp5g3vL8d2k2sfBjPzW7
SPNzaimfMG3iwqlzAoBRjF/HvITUv1T8uTHW+DmC41njvXyaLWPGuRbaXF7n56akXHFEX3lGlj2v
v6aT6zrcS82v27zofBq+zAegK13RwzFVIBaUbDsOJjffT9N79+A/GL5vm7HUMbLS5G4dLXp/SvYy
c9afvipohiJsCgJ74ssq4KfD7DIrzAeAD/F4dUKKj+sBnIoD6bAxHL77rZGED3Pk9exeiU2nilCZ
hHR87K6q39q0YyDX6VWPH0m+Y5+R3xRk+o2F05u6UNzDceEvQpJmdNGCO51W4UT0NeqLp9BzzeaU
fiuXU8YyzANjoH8fP/YHgiJkDcaoAWvpZVd2fSyN1nHwB3rE/kN7fUIXQy/ovTbT6rXnAJQHBjBU
ypNmmSsxBF6581DDeJLVbPWZSnbn9qzj/ATS7w/qEEDuGVV2J7dstClA3OCHnC1ruvPcyTxIfcW/
Tsbw4VD+SZr6GRR4Th4rxDyKRW72plt+MGyntE1LEH/+/1xbOT1dgpDYy+Tn4R4LtRwPoN/CfjC6
nlWczFAkfcgZutxZdl7iouwMVwEpmT1exzyMz/olbZKQ531fRo1dpZXGcaAStSaXouIu0aLeSGzT
ZW9DGui5hT/RR2j35KJpW3VRDksF8wslqvnzqNJCYND1X5pB1+quLS/YKiCpTN4SZj/RYh/EjX8A
cu1Mh24dUPo0DKeHC1yXfD6IZIcHBHxWgRbqvSoTfdu91d1xBhZ/h9FD2Sdsm60SETuth+QsunOc
mlwr5h/Ih5m+XtHitmv4YoOBBl+3mdEHG33EUrLtNcROWll/MrmsdRCo7cYDBwcprX3YgG184X07
0QFXjJtWLxJ5qgsDbGEjNt0Bncusk7p1ZdQYWic5oEq7sn87Lxm01bGl6wXBHJUgO4sMsb3mQLWI
sQQ2IQ8mxlIfeyExxH43plrBu3DVZDqQWCe6ECJdvQBINU8IeeFpG3/MN5fiJagR7qxIUIpt0XJQ
mDsJXIAxDTA+a9a2D8lRl3g2UicPC+GtdKy1t5vfYwuYUw0bJAmSgMFiu/l7ZYiY50zNr9dHwZHE
eT50TTwq0CFCKcYoKhCxiFjlr1MjuxfK0O11mSHq+vO0WhU5ucBQ5zJyao92SPI4IyhTPei/Ku3H
J6wHeHAhcWcRmbaemxMIMj4HkulC8vxWqlI1KxpfZA9VOyOHP37u3rNQzcc+Qrqd0QUMnwAkAH75
RdtDryhb834uc1muS0aZuEysfqoIqjZJYb9hIIXKFXxMvrpUaGs71RYQj07sTMd3y47hAU8zHly4
B+qYQ1SRWy2LN/8thgCt5tIQ0PmZfkZN+4VPUv+y5gWAmbrtgugIdRWoCBtX6x2PCS7YEoPHIyl8
9jzi4rK54bjV2rZ9QydYAAgelN/gVruGXFbBI8ec9syGYZNmotXAGhvak9txmF05PHTMDxo5MtD4
4GDLnbiCYFE0arDkMljb8ORSYDFC308HYjyZBfE6UZ1wfrMQ1V9PfjXPfzPs+6/BQaUySRCmJYoa
BzhK4T92wqPnPLdOeeE82kHtHDrVJuxPZhIIGoWfm3S6wQafNqOEq5Ejxtc29/VcNE87/wyGTdaM
oIvPEG5r1EyNeyYjp5op+CcOsObWLwcXvgG7JUq1QKCjRwC2tsBrW7guwNIklk84p+gG08z/AEVO
I6Dge8PXru9S3oHxKw2ITapokWlFPNvxG7+vc4aMYssaGLI3w42xkOeJDuLMhEk+uNnDP1N03pm2
auGP3qoQ15P7PVx5A0E8W7OEHvqeEywZGn6YdH+yeogmbzSiPrzrrN/0O6laTn43P9d9OmBzRwqk
+sTYHjfu+nsTH88cedkC5EDcTSElzMNJgd6RrXpeEAPQ7EF/8+p9TjP40CyOHpuDMqLVz0cVgr3r
7WGpBWlQvU9ROcV0DfmixlJLw654bCgYeUehILyfjrThUIRWCefQzMBVUoSLGNRQEtQINTlV2drl
J3SNNJ7p5WrB9vb9DnwZy6b8gr1n7hFOPiFnhQ5ELPO/gJ3vNC99r3Xq/Jejnoip5MLKkTh/mRaa
HMnK0jipQG25xeZDvsqAjAkHwq8G+El7tBesJ+u/yaJAHXCrk1s68s/R70dsmSoUnlK1T350Qb0x
jHNuB8OHRED0b9eXV0+wBYalm7qMyRC5H5ydu0+6nI+dOIzu+nvnn3VRA2m1DkgEZwQhK5mwv3zG
pJszTeU8hfonjyj1RxIn+n9en9Azzho6CpW2v5U9DKzes8AYf2M7RacMjCufJVieQTQCONspKr1M
y+QcWx6vvR2JraikwyNEhbI7AMFyTIwc0tF37fFktq7XL69X6rqGAWcAmSFFSlvTD8nax0xgOLpX
bO1ZwE0fzG/pFaSHk0XX+1AAr6XsCc9i1Wh+++qCH3wRHLC3XlsdROFGIUyariGge5O/EgeE6g9n
YQ1CsRgn0vDEkmDDfNGPKa8g2vvnxZsOVyD0QVhmTZU4bWaeNwwIhc/bTytLFCXtO0VSxW3TlbMa
1EJtunh2NUMj7YB8/wbokcxzM84aIjbAZTjRVCuosvL9ILpi6a5VAALa0iH0xgZcgCTD4XdwiFET
f0yMGMJHm2BXNhdz2s/zo11iBEZLZ2tfJB3ahuCGfaZGqt126Mzuk0dw+YLHStBsrAWpCTlrYvxi
B3Xz75wA3Qusa6crnHB2949Y7NfWtu2MjmcA+8lsZAhEV4fML+KKyMyYYcQv6KfM72FvwpF3U6km
9LZjdAD0fsa6sl5Cy8KBHuYhqO7kDBBzDTYkTBf21LIrdykK0zayeUgMCuy6IFk1DmmDngnQD45M
9D4XItcAPgNa2DWT8BBS/fsvBUo/uOPFNcOEVzfRbcelxS3PPWWaD0Uz69B1ANkqHL6lgciorV0M
HzgtWhb/epBD7D4Mc7qR7Q6zoj8k5v2ogBtgcdgMaBOoirU1Tzo1t2cs64J9cSWWH1HhU4NMJe9Q
CDLdhN5+ZwhmySLKj4DwE6bRJBVvStcGyoURjnerKtJzn5m2Jt2y9F70FgVm1HfHs0kMGCqgl/PF
OLheL5kGCSO7099x+FBzIO0G28Elw8RsiPWHODBNOpXmYOwiNp2DnnK6ZHPZWH9vnmI63QzTYYgt
uN+BJ6O9bP3oL9Sw2sEW/oSqd6+N+2WKc+elrOK1/ZdisHhFAj6LK6hlP794LIJW3R1BAFCLW5t+
AtF1dDfPZGw2CUqQVJa+m3gcwHedq6bJIa963M374/VwUwa5QHOpJbs9y8aB/pu2/9x1N+Q8D/v9
sp2a6LIYC8SWlAYAd9XTTKUdozVb8joTu7m2kZljMFE6OXg5oviRZdmrBGP80nqyC0XYU0iLT+OZ
/9EgRy1j/dRf3tWTyQVmUAHYKeYzhj3c9DRNURuMqlnjwVqsl80H8ZIj0GtPaUFY7izL4Eegc4DP
nOdxcAxVKLpdsyKC0yMhjJeCUhopXO8QqToaGDPGKUYL7IQ3DMqNl1rNlUowhSeX7FJ4DiKxP/dO
pHv5Ppt3gmRT/LuzsoqT2Klg71/Fg9BcCYS6CKsdwbMVdxHYVdp5+0amDfi8oSvySfK1LCLECQLl
YwPgfB5T+mV9jtRNCBFvPeyRdmUpUPd+lRjljO9eqnUcHmLrQi4iF0XjWkwQgDZqaY42A+K4uJ1k
/gl9K/kLjQH/UvHCTO9laInFyseHO78v2XGX6ywcKNy8Hfh0RYez1r7qoQAeT1GVvogOsW3qAPNO
Grizt9Z0HNfKC/GH4T2nett+M3HxOTsP0n9REQJSTtIJQjv4JxDfhwq+8pnRj53EYLb5NXT4o7we
37sQ0hDsdZLlOlOXPAt5tFjL7fjSCvfLwJfhom3yihuBmv1y3oL2owgyWCaod5Z7LmFy+SFIf3Vv
qFzxGkit/v54X77d6mMgvQX2T6c7xnGrTRsoGQOaHjTqfdZkLYpbzdJiovIjzgyruxwyXSi3UEf8
HbM//0zNhEyQ3sB5mTJIlNlvcX/ADLetf5E9eXF6yE3yq/uTV1YqmVxmZmRRrrfYXibJmdahwJKg
/vhEe4TfkcM1CD94l6X6FtZtgmv+aGMXhGzWxJmIjwYaNAW0fWi/L/GXczvdQSmukBC3ZmTLsyEs
1A9Adjga7m0oqYdc1fQDK5b7uuIGz9yHpInZvzaxY93dJR8ukS8KAzgiAwYN2hvXVFm1/Z3xPPZC
8SyJ9RM+N7jI4giL2Y70aAaIf34kgk9EQhCUyrv5Yr3wHfK/8A4BZlcj8ACaMx5tIDeCJF01urE6
NkF2W8TKOmQ5H4c/S+pqmEACfvEByD7Bj2LpHu4iv4f3/fybCuMw3ykZGvlsTkL9ZUuVdrVgAQhZ
enZiBI0ryLjpu6cRnbZ8c8dWuQqBrkdFslmW83pK2pZffhQjcmpC2uMS/5khS3n+ktLbHnsWbnTC
cCyZt7khvs30WLAwCYN02hwXgd9cciBkbFTYREj7AZiWEOsfkXm4aJ6KvdRvxR+FMk7koddEfwVV
eosjeLDk0A54W7TBNvp2RvHP9Kbmu6lcR4t/q2iUMfmO0Wrw7HJIe4/bt5uNe/Izl6UQBlxZ2k3c
Jhvc9d59mNehq+kPka0KQ4NnT8uwtDfExePEzizgthxzjeH/TtlzEhzbcYv0BnY+lRbcQ1Dtn8Kd
yMbVOKrF0xPRUnhOu8ep2nt/+DVGQYOLW9mo/NI73HFEjXMExfoDhRqVwaUoXKUknZ7DDSrJcmAg
GlceXQDK8WV1rV1w1rB/wbAGEZ/J8Aln2XsxM8wop8sVWdX1WQMNC24tQwGGh0M8BvN2R0A6iyB8
Hz4UavjGMW+VCvruoNtm+0Qr1gY+WLKsxjNFW71BNCnj6NdTOVWiKbTrwaJaZdNVXzsSCrtd4frn
EKBsOSomExjpGlrr23NRTRwdzMrdkZtAXQRO9EwCIvz5jakpNu0Te6tIGIrtYVJ0HamKx9dzYE+6
JOWjOsy3F41KamB2xoMv02M7TUwZKjrO18T3D+KCtTN8VYw7gMkihQsbpj1Xzxydkm+H3jOaAmYN
WinUS25SfTq9suCI+oRmlRAQDZJYdK3SDZaac+I0FXERGEMiOfhrzEXCt/zW734Qm+1S941Ek77w
xq1pMXrpXUOhMhBnzQ0H+GLJuxAbC68+N7Ou1NBRbtYtbAnuK6qdgsKkd0zqDyFr9JWSDpBwef7k
n5hgh+BO9WXhnlKyvAa34StyXbzN4tXau7e26JBfHRhdEAkdv83Kqt8YHsVR3nvkDB6xTqA2K3rr
lA4/Dabq2A9w7oszoEemXmUTmKU1BpCx4zOPAhDiTvmamBozoKOyzloJbJg6WLegbmguQgpddE8W
Uag9N4WgaTxcmYHd6TUoAkfmxI4Kb5YC56v7A2NyDDmpcxp168f2surU0y9xlmeKt2ZGIGpxQBZV
eg3XqHRgqokwpXsnHipud+RyCaK6/WRqMLwoq9JsmG2Qd1Nt4AZxCUhalLpRIsfNEOdY3BY9mgf7
DB2A5fCr3zaJDy4SFCeCB31qtCNh1yPysdZ6YuUkKMMFUI5vBhAZeKU1AhMJP+fW1PXW+JlfzL5T
bFqPAWK/rCEp+ZiMpl0X02hMFhTYdnAuLjXsMOt8wILhtAl0hcxY6n3KN8XvicMh5a9FjoIkz++o
NZW6ySIY/ba3QO/RfxXwPm2zrK5yKsoEcQN/L84F5X/wef6vF7rEXoNHf72cnNKpk0eRB1tlAo5X
5Y8p01iGykNJE9x2wAUnHGKiD+NiJuzxVps2gOKecZXHFdbffyrYBIIn1brOUvnPEXDA/8y7aUkV
hnu2hcoqk2Jvir41RAgjReMWgnM0+meSina6gfS853s3F7PYbYCLwzf0fW5Kpmp1QoTrwNFvQVBT
QHkxEuLOSZzOeoJXNlYQ3DwqVRSVnUtfyL86vagzIVlUH4LXrhiX8uVcX2A/GzywU7p/LLo3QDGW
w5iUvFjr0EAasXoPT68cmLXST8+TomSNY830LYn2yEzBokwbi8/hyLUwa7qxF3ynNqZaLAXfs3w7
xpZfhwk1i5ni974+henr190xEljfK4YkG/8CLcHePvJTjxmO1/+ZiMXlv0G4Ecw09D/CVgjEH2kr
gju9Ath//hgbLR2KjZHL/zO6PW8lk2d8aSrxGeF4P82nx+wjDbgMABPZ3L1FMVOf4lFpN7E640k0
yExL/5HfIA7XuCHJgUAInRSuWmu3qUPAYRFRiSwGuhtdG1duCXGLavNjA9KxRzWghvD1kCeneoOq
HWCyaZx4j6IYe4VsaCbkokSYcFq7yV6p8mzrtI3Lc/XD6/mRh5D/9sUlonVa2JeKPAkw9NKV/LXy
+tmRz/vCzziDjwDZHLXLw/7TRPLn7PCi5/V8/5NiIOHjIq+vq46TrP7SlMgUSnn7opjOUcDTRGyH
yeuZR/v+qPafl6KYjQvyc5eaU6LfHdnwHO3u39pZnSVyIDOe6mrCNJZqag/8uM0ae2yUv3/6m6e3
cMyPNGGkl+5FSNBsq7Qa0dtOeJXVgrEgcXJyUcnc8H3Q/6kJivxCgbrUvID4qHu86GErAZLZ3oYb
zcccgZTP3Qc/gLKfTV9h3/tRlCEh7bnjl9WiTSeB1HcYSAUjNw3Y1aiAnVYDdybvbt4vKQuQjlsI
ajcDFz51Eaw6vYvvPrF/+t5JDF739sdfHWUjOe2Cw7nNaUbTbImrSUtX+q+d+TQPqPSTY7fSmwWi
JBiB8xvBcYV0oPmKIoB6EF6dt+nfgLCQm+/dEW0r/YTsjLrs2tBwFJwo/gyK8eYBTwk2q/iqyiGR
EKoTIyQCdpovQk2WQLDeWLSxkiCybvkZoFTXSC0Vhl2wqrmqHTHWCZJ6vw/HdeO4bIIg7RqwQGE3
ncbxLMiwfg48EVtrh7zqE1Mif+9U71mrz9QJ3blJCOm+zCjuIzNvPLYFoXHoVb/0iGJGzo3ozkKY
X66zo3iY03FPT6TcrPN31VVCAUYmTEAGzp52oecNRd6lFj53yOo1iXTM+1sm+XFOmZ7ResW5xtgi
mGMCXyM/AvY7BCrPOo2XPU/lFGpo6UW+RXAHm28GNVL3mFHN7tYyOd8S8cuppsHnJ2hHv930JejZ
wCNdZpJ8467QOejAcxxACMcJgFIYn+peAuD6/uHF8gcfMRd1Iqpy9m8H8A+//SIqKAF6WdZvvrAr
wSXVypBsnii53nOMIeKUiqWNnJwIpc2cQzybx9zUQRPeNZCLV82/Xu1gbu7CHB/Xp10tvajva1CQ
0LlpuMFSZ3+wxTBfvuMUI/OkBXXp4k2gt2bct/odFbzbeIM7UI4TdZpC2NWBO8rZ7AzVAAJQdtro
z9iXArWnPvliFImYThyvPnns/66bHAxN0Zg8lbWwPZwEcYrOMTbY4BQZNsxJbsj9TBEhr53CMy9k
LFyIsZi8GC9BXB3ivOujHYeil6eLBK4rpuJgEdiEfB84F5O3B8mxk+S2l2nG8/pIGnJf8ozUP+DJ
PbN6pDRygiqke0V9imdhm2RaqAQc71tgdX31cqOuabkqqOtbpMhAXyTO35uaqn10j906sUX0EtVf
P346EFiTps9ekI0BadlVOa2j/whkfP2udI7Q+38umLZnavNVYAshTMfXlQyaiLs+LbAmzh66fiM/
gHAUxT9SQ4SVRkUSw1a7RFnlQLrcYLxjOZjqxpDYpo53ndoPmV7v/fP8wL1IF/S5N5/29xADQoex
U2SkXbVenXbfn199JCEoTwKB/qqky3pdNZQ/mLheSYaRkObOBvLqE9TP8HSh67qn7HYbudHeA1nx
j0CQH0Hlr2qRR/XxnAduUF6KPYNXlHwSkqECfp9xFjXx7UFNw0pKoELu9Ju7a793PKcd7QOMs/01
5tU6PPevVBrYITp6gj/GqfMUPSi2A9F98N+ohm5nvIAMbFbeE+spNAtDVSVAzgt1YsSJafi/fpFL
HlAf/d2+IoqlcWFTaYySiLOH3S8vJ7wYVOeu6hBaRdkT1SpVzIn3omuwfkiIojLuGY8B1AS4ZFV3
zD1DbBl+nYa+TuWbTcKJlke75qP2r/bj+SLJSDsd2c6k/tDun9hBsNZaWpkJeqciATcqAvEV+Nb7
kTEAa1qEOT2eUz4/9IF+bSefRRGHpXWAxFqa38RaDZ//9k+l/fsHvtqsWV7+nPdmzx3msFe2ItLt
U4aKtdfB81Qo6EzsYgJXd/r0n9WM4Rq17Wn/yuE08ACxzeVWEEzQ+kUIxHzSAIXSveWZi2QNNft8
lAJdANtl1SQNH8Su1BEBY5H5n+mHjAf//FXNXYVuIcWtAmDn2Pzd3iUgjcxB1ofAIbqaMvci7WEF
zUXcB9ciofpW3/LRSCStbyYzbRCxHFbHOdHFGOi/gj3xxG5YkioLETGqg/0zTXsCuJywueb5TBXS
7myiuWoMNQrtSTX79A88oQ/kvt4cukkPTJ2WK+6o6CeWMVJpKsHdD4V7cuyHSjTYmaxj60A/ihoP
rQr0fDiDz/PUyDkymwKc69TBpKh8SfjRvVTVqt5jtQ1/BkPGYHQlzcgC/kKiVCSX8Awt7vexNLRg
qZW32lIqBtlTBC6Yghb6zTiLd8QpwfzbmIFcGcylQbSD9nFzNVYE0ZmoArARxvG+m7wn6W8gWuW5
a6affpyxs9MbKiqVpzPGZJvSj+3qUsVzLkg6mGstlfAx1mXNlMdTKWj10dRo/nFWqh5upjCee5EL
PkVJA1o8FMxtAPTqj//AUlK2OlI56qtQi5qCaxylPFrMf7A35v50ftsblgTjyen4h+4BuO9Q2tGi
Tuq8Hr9jPvUa8ZU7B17XvXV0dTqE6/BwBYWcQDhO50DYXaBU82D9mZpbEfK+5nN548SXD4UivKCw
plROD9rYO2mmTQCddaNsNpsp7Wz4uCpH3vA+6Rfkclkvg0MNqCQRKYONZXIuVlNC7HmfpJpRXeDd
/NZEzyg8eXlywF/5NreFcUUXeHN9OebdtF+bLqxEhw84zftKlCPTcv/ZB1K6VLt0bq86FwmWqj9A
Qi4nV4FD52BLL14AVCEtTxMG50+WATVOgaLpPV7NRmweOODUlypjW8xS7gveuLPE+QcwUxqK6NOr
Zt1IPR+0JqfZ1o+Fa9NOW4aBdhVQ5cQlss6B9CXoSqmU1hrOGJSuQs65jzqxeoZnGDMSEGeo7dAk
d/xovX/hbPpSIWwBHoSZ8FFgJ/Yuz4v7J1UcSOP4n3VBw7DZQkEXIfRUGMPFG0Zzr7ml9U1D2etA
55kOIfynzFvEBCwUU6zm0QHTxdjnwECXXffXsn9yYw3N9pQ9ZaHIsdV7Vw63KWw0OMCb4ULKzhZ7
gKB4JnKL7aFy448+441J/ag6J60dILnBZZz/lKuF+IG5iDhqvEh1dzyWQp9VNbBZCgT7NI8wAL/M
N+3CcHZH1m+brO0OszHTdxyhPjNle4nkOizDzAsIMgtKEdUGvpCvmHznA/gu3iJHfFb5Gq1mtkHl
6OS6Nt5Mpg2nPuAJhuj4WgQw2TmQlCv2xERx5heC0L9RV9Hi5EpDRoDodt5VuT1nPeRpL1tdr64O
ISVg9Oec9S9GUwfAPmSVrD2vEvjfoOsu+16vW/UqZh7Mdcseyjtz0i1E1JgrIAriyPwt86nNb+mm
FbbiEd/GSybAiZWpG2B5SMe5kvRgeYT2vxk6ijPVwnBVUfTeZC1Q50AE4YTaU3TXTSar0yX3c3Um
4YUneLsqOcu2+Tk6Y/KG+xxl8IbUCs7frq3usUyi7tk7RpEWhboGRn4B2tMs5IXmR1hMSdTKd2UG
iaag8MMcuSw4+rxxWGnCU/wXU015N2y2PHhTen8AzB3n7JTWxdSOfVPIEdhql2VB9g2ZxCet+VEi
kHtq3G2AApBAh7psDtPPL+Dcv4UMNq8kEbASVNn6PecYvYsGGTjThx+1LdLvslbfuqnlAgneTGeg
Gu9CWQZEFzrHhHcI4+sbLwS3cpZMeG8OinfhRoV+TXD2Xm4selRF3XeGa254rsHC4cFVXDjYDeaF
55uqp+Iuzx6aY3M9DTcRgsGJblGkiu8MiT85kSJHwSkGS3fM+NKuhZX3eYhwaIxAnov/RDC/4fhW
Nlv2VFiDvgKm1Uk8w716+XLDrqzgFKteD0sfThQ91OQXVvKj/+4QMHn5dxCtCaKPaIqu14/hhaW/
1Mkvu8ysJknZKF8hVe7U6XHgZAKeFxXb4orIoQp9xXKyRiQPsE9VZ10jyXTJ5jhjHeFK3LHlWZbM
DojttQqmErHxXVAfmAo44OVtGa7zI6yeub9mN5idpQfzcsliOXL62ZAZSrLescrnetm1IA4oGGro
jSQb7WeIyaCx7n6ziQa6v82BhxtZV6PKBD7wJpBDqZDL3R5pJNAdKO/KSEom5aSi6rYpD+77J/bl
5XezuaNoOpE2jvqh5RxGQCNw8HcFd4LNR7UMaRtMorHzfzqRxHrfmEpXSRyx460LTA9K+EfpIypw
VrEkSmamtyQVIBlGlGKGVcwyTVzwbIoedHX6d1hfd89wucBFinP5NS+lZmHSXZ353ZLDLnYQgmuL
0B/c8aGGYfp5srpNnAoaOZDW6Y/+jQDgLUQlQWq14mgRaWRqbQxlN+r26RIwNTvq1D04P/gLrumn
0QXs1rF9dxMqABzqTY9n2YkYTIXTSq9GOTTDTw3frd2+T2G7FnEtL0m6v4wWapn0ROlxnHU6OSta
J6n1/NCbXziorRmsdSQI3LTjQqc6GSgFC7gXL29FG8+/cv/tRGZzJK03+BoGEKWw312Vl8AC5Aag
gl9kzHNI8vqMeN18OKMujVD7s/7CR2UKcAGDelwzXJID3dovWLaMFj8ysb6EyhIIRn+p08eBEWXO
XFsnJPP8uZ0fp5R07jcnnxBLskkMyVmlB1M+Xp0aNGndizGqgoU2gMKSOvRJHv6qGL9kbOwMjG27
rFTRyV1IFCwVMgtdj3QNg8P2uwFgpNHdGMra87UqRlyZ4O43BvILSGGIM5CZSbLmzaXl3WjzfhPh
+3Z+zYb0l4H81gPNIcJ8W4bXi91bq5e3P+PcBeY4ehGR38bliekuCDd0UnS5Gt00FQ4OJ602Xx9M
KqLQWGFcamU3lM7qXwx3tBW2SNcRRRLaCxqHT3yKIl6URkKXjrptpQIfnco2BNKsFbcE/Ncz0+q2
8GwuxKIJoSaYN3h+b6JQ0HXe1eBrw+UC9ZKkwERPdPRr9l90+wYuJ/NVZjnHQd4Y7gyig6ctY3ac
Wjf+vnZyNdO/wHKmiAMagIkurc+haMlomTjPtyWf+D22FiyhAvD+gqrgHA0QcLhXXcPwk8Jj2MfT
3dD97R23JMMTsOP7gylO0ekEdffWl1NvFsmXh51t+yt8AaNjJya7rfnlIKDeNJnf1VqBiLiJo6tD
uKDcT4yR3FNwMBp2AaJmQgjL7GCgksjoYcjn8jbotX8z8O/irNjIBn0l6CcLF+L1nlPH7JS18/IM
nY8H40QcjI+h3xdHeF7ShoqL88IU5S4kRiKonli1T+AuMB6wXoA9Q6T5jPE0sF6yYPP3C2D9lSGo
sYrUDRxphMSfpctrgmfdNUmYv1B+1tNhtBl25Frm3pdmxqgVf/qtyGulIkV0XlBY1QztNNo+e7sA
hiudSyZfEvMFenUp/FtoxvQbRUdKVVjd2GLOXrtfBZDEwX7lOPFU3CmXj0Qh4RcaOxCZK0XMvL5k
N3J/LMf86/0He1BArCLzlLHFVxT1SI8WcpISio182blTfbwf0ekHYS8b/qmmMessT5KEnEna+SCl
9WcxvovhydE4LuvVqW0KrB9IHhCvlREHpWXoh9c1jtf7wgias2xMap0ufSuRZy/+MahYX5ads6OO
SJ6ChqMMUC4jaIJ0axM7h5ZV/wFrkYipN33jWAcgDG2uUoR+C3impt3Co/asTSWT+1rf9OFm53wG
4DePb25Dx/SHgr5TlgA6kmlgQ5UV05NrvN8at0b/ZY49OnOgfIhPnKDu1c3ZHePlqyh+RdD4isuM
BhmCfIut6VvSJ1lVMutKkSXhzk61z3bQAFADFX6/ghXt5Z8d7V4J1Wsj1BuavsOtGXy4pIYZC2Az
TnULvexjCJrsD1ID0ky0iebC402EgUwuZTxqrXy5JcCV1zGptr2dHS1TMe7sBwx/JI2RJDx15SXB
r348WtL1TllGXiVxgNQ4crRD67Ocv0s+8/VrRQphwwhFn0yovZaEKIJrMRTEd479B0fuJCs9jrdx
dZlh5QOH2Gk3jg6JhB8FUldw0GHzfcKObXVybENokAy/Z0JZh9griw1yPRu0fPqgxdf9aLspsUYT
U5uQR3EUXM93bdDgTfFp6mCDBaP89UD4cWfoWuKWHS/1iBwKrQwl02/wnyUV7lDiUwGKQdzG8B7S
rjZG6y725pHXpHLR8c4twSBOzg2sjx2qQzYyFZKtP9abKqACGk7lu+P5qeJqSX3F/4sgiluCM23J
qv0C/hxLXEp/xJ8B3Y5eZAaBEoVscoXCnOAEJnaY3LIAMNYAG07Cg9QUw/xdMHX0XvZ/daA8f+DA
kGuMSGsVkL9YwcxmgeHTTAxAmHiUjv7wFJGOMsIXPhpGsMFN/ne41teFYz855qnLihGvOTBrQX/r
R7IZZLQlkUBqaaYWbyb22a0kSRXJcjgmvrHBx1VRu4bZ7F4Wh7RNMIUbtBLZXCfosbL4r/x7d6Cf
+s/aQ1ZrSYU3tLedK+vIFH8Tj3jTB6Xy7E1lxTLrR6Yveb7I5FOBnIH12O+jnVPw4BRfdA7K1mSV
8mccahOKcAcv2Esm905CFyM0Ml4CcmPvO23CnstPjaAFqHE51DHXbkBixTkyChEGjzOWAkRreLRl
Q8WEteJRHSvT+iDTKMKaM6vqFjZuXtb8P0Xn+7dEVjZ+sDoK6iV35WULBFOFHvM7xWz0hmwogEsb
fnBUqei2nl6ZLx43ElKy5flAxBeeP2afhVCfQjiv7EXc96ahhnrVFN2b9Z024pFgeRsgfrREd9qj
SPFW8ugDP4vtnXrLg0rh5CYzmHouaGKLFa4f+rffY67hwpBykSVMLwleg7KbIClXyXuiyWti2wpx
lD/MAx6o+162/USyInFSbQ0d2T/mo5G0/UMzoa9Y8TlOJu0s7p/1lFHFFQERb2/V7HnIAqSPagiM
MAMf1w5FwPaGNCOcqzY6ui5KGucfOdqIdsQsL4JomcR+qxTCi+2jgWUEEIWtKAlnHlW1nqfsoHYC
53C381CBilD1wYwwZr3Av7DLIYWu1g9+1jPp8ABhprGgRmX4+aBQqYLXeGFDFmjFpYMB6W0ByRR3
lLH3otijFl94VTzzkPG7uq3jZOZGK4CHOFUgnRM0ZsfRBi+VFweut6J4ScY+lpqZW/ZDlzwEZSyc
NVcXEj3lan6U2tooBA2BqK6sFGonbog1Ak3oYuhuDpY5YvT64HdlOmSrgJrg9b92d7AHBUuzepP9
ugrO/q0Zocdy4E8u/RicrzUdizHGSglaxMiMbhaD+aPCSZF/CjsvmYpwVIlLNtGTUDOHlZHmTKoK
pl02l+Np7XfRWZDuGh0/Jew0G1IiJdmnWvnoJxxt+luWuHcFMoVSDrJ33PugdCSZYN4CYyZha7fe
/Af4fagwxHCPHl1VopuQ+e7bv0tPGKxdZekRqGrlC82peQtinGbjNBX+CH2pOJ86xI2oS09we9g1
Gc8na/QvlMtwxp8vaOjnaGA6AoJkLTKcRLi8tvMULPRJ3wQhAm5Lq517/dN0WJQ/Pmw6cIU2QxXu
fK0qxWbXEIclvE3CZijO7l4S3k9ApERvHwFLppdedLFwt/M5VO1ynMlO/P9YEjJMww01hyMuVRAa
CZWxTVYiBuX63RLK+4w+3bUTd1ZTbQWxBG9oFj+oW3ajoh8+wBh4NuKQCrMgWuCoPYQf2ILa09DF
lBkssYtDKwmGHhSxXJv5mMCGLVsGOMR+TSIclOB5TYrd+5P2O4dh10XhF8jvf9iXPluf3bYTAmT2
Cx3YbiO8jTF08pBxqOgPY2ggN/FwLQJVdf0HrurAma3Tey81ufh1IFsqPsBKHq84KcYE5hNbqAcq
VJCk5wV+jRjohZEewF4NaO35yptphE3Ad0OcFhpbbJ6d+EkC0G8U25H8lS9QzjfNSj99TNM/r7Kg
GuWSmISPsVjyL30UKMXzle+m512zpBStDuuj4+wtrRQS4dkeb8IH3Al5Ht7bONzTcdmsxvouvz7j
oO0wMEanJNkoMSglZCtPyFwxRV4G+AOp3VazPRHpvIlL0EQ02YPWeohukW2EncDCk8kHFRsNEchX
c6jJjTiQhJA/0esPOeVrOPW9Pzn+wHOGHFxncirK2n6m47wN6Wm8PQ+9wrfJCRdP22nBUl3H6Wd5
2UgI5OnCDrFHOZHQgbe2iOCHF01Bw4rZI7NgmzbKG7IUYuBatPvRd5rCclxG3AoT4ewFdBvkawet
eL0DR2VbpeeR4M6+G1vejTI7nKE5c7r1N44yK8gxv2167z1PLmIE9X2P/6E0u7utTtZAfyKDjokF
xsJG7DhuAul975E2LqHuts5Kai9uIGxzblnvnX5Ji2aPhagzFEkh7MD3RfNdqGN+ejB0/rSwd2/g
fXSIfTtuHPQG5FqUWExMjY8vhDGrgBQFIU9FGmFXEO9ruh+GnsYb1XJMTUJw+hZ0iqYz+CcE6fmD
QArPdXUH1mvbV97q08O1zszM31kGUK9Xe9txZqH7p3R0WpJIRsjZm4K8+X5592wGWCZoP2H10vFG
dWr3MvExsesqAameAPw692uSUmctCoCTKOPlgWKHo6azmJArkDj1LUbARTNzvtbK/X2QT6M1Z26J
iqDLH86cPwVrJSEqKlFB2rob/aX09GAd91znnDWLLtZgzd99nPyKT2hXsQ9z9naH6WP0bobsIDTm
ZMavi0i6GrlvuLxaYFXlkn1g1ZPQstAbT/H2qLNdKntFyecqlsxy38l+Wb8glcN8j3m+yDCAyxBf
9ehhPRfTKZjc0At70GcGTlcodgVvSkijp7XkLKVWwnnbdI+U4NWbzafda1B5CLBHmMJs1gwahU7R
lL2HRS8daJY9D1okbkp6tuC3ZMCv2HFirifqEjV0lPppLRAMPk7aEj35qz+tL2wnXoUHeX3tTG/r
oXeAzVX5fKHQs9NC3wdSH/olQQPukrurxSpPvjMyPucqvEoZs37ElrR9/iTfEOiz3lxlcVmpkO7g
iFpTOZKelyEjP+uHiXmXmcIAuo4t48clZMy4tBlIrn+HzxtrlLVHPiIkSfNBIZYg2vl0qNFWO0Cs
Z1pfAUOMD3XH4flR1e1CYEgTFTCYYV9UU34WbGwVMkT4OAqFCdAaWvd5Zl8IPKJep6UYTRFlIyQP
PfK1RbiwfD2KB93MuFaVmFh7ZQOq8hhNQ89TMSdwTGgNs5yLfuhEbhRQxMk93vCbHaBuFLpLc/NS
lEbtIud6Z5bgt/Sz4ALMFJ6OWoY604TfGXlVMabYGUPOZtzCTb9XD82GJrj8WVE+4ENGoCkTxK7g
yvnJEz4KGUkVpO4UpovyMRH0peLXMMqiK5DTKreuDdtrfz25NbmOGQ6hAQScY8vI7U2lA1dwoupV
k3Iop5T0CBRX0qkr5vKKJcw4YA56VXm2klHsm18xOxPiXpNrh8uO2gnPgp8uLwI3V6KLT/Y23RRQ
NUERlgladnFZzKqq6vnG4SeNQdYnmM0BBW3i33fBT6vKCDcO9uaBCll67PC/Xl5IEaxlOPNqBQqJ
XNu/th9xtNR2uiJIWgSbYt7RnEiKTPMuU/AIheG3sxdHoSljraYqpVtmEH+kfuhSbMtbx+mdkwq2
dlvk7WJ12czVo7vTv0sH581ziNFoBv3rnq2BJMCnQOinE+SZ6KyXTrWLITPMobVx22H5oF6iDW+b
HiGOeAEwfQe7rqW9FR8+zWc2WQ8i3fG5I7h1VLacU6cvqUUI7WfEWX6fXi2fGZbhx+cBPvUG9V8F
eLiJVfsxEY74QxyqIl6Qbsy1teGBpRsYUUYojnj4VPcNGSqmuF9KpJKF4Su1+Jvjr/GccQ2BeuTi
6ADC46TWp/1i2lRgy3LBK0Nent0V0hQdY1iH+kal/CScSfd1lQgDep7UMWHDHT79h1Rubbiz3ijA
hnaU50NPBYH3usI2w/UGcBGh13Ifdu4PAM+0SmDkCkfWVNklEmLoywZ6xNiO6qcXFVKX9clYdN7E
7NAONB8B8qmeCUvu3SG24M38cNJGPcugnHxobOzZjbfZR1X6f2uT7DMsp3maPRQTePJNR6r8i4Ta
KFUoxUeKaGW1prOCzfF4yzk1ys11pBknuQcC3+GLpx73TUZenmDgnsAH83GrWGpWnyCY19p9L8fi
lfg6z7I3j9PrKznSsZecp4R+MVHtPZAUkAABWodwLgxHwUrGUQaecEK28AQZbnnVoA74DA8rBxm2
ZGgak7+iK0HBSASbPyPR/hvCsrKlrrgOtaQNh15JHWv3Rs2XE9ZkPc5RMMMl1ij9XkZ7DhGmcywx
r72eK0Gy8rohGWlRrjRt8vFM1jo4xRwbVduE9F8PE8PSqfQa7GAMP/q2I/ibJcTtqlkEsandBtiH
ZJGzuNxn0Ti8+zqjyxSpifmaXR+fc7lP78TVO4+4UjNpdJOA1zt+pU9aCAKKm8rZ2+AHcpG8v4xs
9V63NpXL58UsU0ohRuJrEDUsEB/JqfgWHeu32X2Wi/aMKYMBDw8RQvgpG+wWIEN3ZNgpb/5aXeQo
iCSi9G8rrSnSG/d9XcruaxGZck15GIYpXS/99oBH85UbguyPafto9l3ka0TNpfLio3WX/5uGnmg4
sLCn6oyqagoU4XaOrIA61DQ5V16ia4utdxc519o7VlbRljlSlg8JnuxBfBYPAdSUpAfxopAMOKxP
c+dgxxFfuSZYXrNMMNkmoJO8CPRYIW9Q+y588tvjeLduLJb4lfFT3RQtxMAEnHj39vyEbg/L51Vc
S+8/Wt0b9pNIQC199kCs74h0J+OQcOr3p6UHEYfS0LOZMUxvZRnp6GwbT9T7hr9Ifa6PJUVTc7xk
2ew8nRb0p3eHBZ5owTbKbZBwHo31rz1WiZhY6W8StFbEfM0V5ypxljhnpZ1d6f8DKUK6RQwFuNpZ
+iX0yyRFpCFkH+CMDptmRqHVOyqrRFsfiseFbg5JEUtWMcaStNxTIp59S4cSl9eSecpKlxFbXHD1
2bywcwDQd1AHZ5kFbKEY/pl/HAkXGSHteZus4V3o4Xib8IWXwXgImdYKbmSxFmOmK/BNRHkpbLmR
LtabRkJcXi5UIThQrKcLtU6WWtmt3lD4WVJoSBFyOy666mqPAnpPhbgsGRsB1BKVv+8585/ZrHPO
KJb/oDkGLgyFYrjHWu0hAGySwcExKG8MIqIwewc4sf7ffkn4o2pveGCF9MUWBTyii/mfYCGxbDsl
d56/0bVQRcJBUbopBx4ft7lDVNVsIDoNHgCPOG5PG4Z+45Ehv8lOOyDTVbm7usSpP5rOnFW4OgJX
TggLsSFzYz+ADYPP0ZFE20oUMjAU4zrnqtIt86mXeib18bfpURYGiKZ4Ho8rGcfI8RM8vt2tNkKo
swoJGIYifWFg9CE5yjVnfXfng70aO4Z0R34zP0XgbOf0ZUrcKj8rtfE7LFSHl48vxPMu1lPreO0A
Rc0g1ecqkXmT+uvjoB4HCfCJQC5OgqbmxXBuf2yWEDGhIDvztJRux/v6D4wqcV3o333s/0cJV6z2
eowQeLeYE8xDNtgvmcV4W1Tc5oMgiQm7ze/TQd0+j8rCH4afrGovs7E5hg5ynvWnOuAw7yjoG7WZ
Y4WUnnagJUdMy9Dcxay3XrEs5qwhQC9LyfkaZAv7rV7f6BkO6GuEu1/TU76yy8yqC/5fG9XAzFyi
OUQNbTrmTnTBWcPO6dtNDEVHY0indSr4d0f2AHrLkAcEJu6FoAmwc7a/dcrGy9Ybz9WYdL2sS6Kl
hGzq7N+Z6B46JKr1aakRPlhxjlMhccGyoJCu1iEX/k7+l2pad6Dq2D9ur3mAkkiPpU6b79X1Z5eK
bkHPl7UOAlN9XeqY+4pBhbZwGajHfxjvMDJJe73cfBnYh5+SzaAkayIs1EzTVrl/1duqEWGrIhG6
1gc7Q1eIXa82IOUKcezMi+Y0DnCnWkb6yf1uBhTjTaBf2aQK8dA20K0d6RbwUBjodzbb5Y7if2Jb
HtpG/D4z8KLSm6AMCVcpUbYUfnS8fKScRX3BmSBhROsuQKJxsyH2rJMa55yOY6YQMRFHakj7NDzk
oBjV6ElygResYnefvWMrkyrkwwbmyI1CQZzf3Lmw81szmYWFv7kj0SJUomrT+sv2qbQ97zQFsxxB
6DgPqQIbm/UsEvhXxx5Ng930TkRXyNxsA9IugwYOQ8AFXkaf0MC1N+aHnBOhQK+KMVjieW3TGYDL
po6t40mmXRl7uWq0r3+Q7Ph+5m16BQmdqdUzhpXDZBPQhCSgo5FVEQlxqmy6VMl8pZkqPd07TV0r
JWLB4uc8t41eryfHz9hgfg/o9rWDgDB16xJ8PymlQScFAQs9VePXQMPV+etKTXBTeyB8k7X3FF5G
L57BKtrYQtK8tTWfdlEBKtSUehTNrQ06YIhlcSWLayrSX4bn5+x4IyGLfhKwFyA+gsSmr5Y35RWE
yW/kabmvGsev5KWSKraROmZNdI3oL3loJPCT1QvNXTvZyxfEmseC18OI8mWYJUrTntvauny9xy8W
ZC+8aslz8FirIgsq9uV0JKzT58ixabSg3slleufa0JVHqytFgw1061a9yORL/FgHskQt69GguZya
V9FkydpznciyaEuouCDEzLdOkjErHoMdG6CJB1u4PXHYJ7c9Tu2w7CbecvuIKFdwlcvAF6VBMkCh
M1mY6bsTAY0DX7PXm0O/FTiQW3rxm+syUIaRa8MUe0+Jl3aF9kg9ifgOkwfppbkttgx0eLRmWip3
egiigRAJ1LQFpUE4rnNWeNuQy5452JMITfWF7JXRV8cgEtU71GtFH/M3UARmlbvJpQMmzpoSUHHb
Hc3AYi/jXFE76LPtVdRHH/sfMb6W3eWqP8X2y0LqeMh4m8AVQqVb/IF78ca7Za7VkEDoteYRYMhH
QmGsofLRw5wwU0iwhSvbWJa6cnf8/CNkj3adXkZnzilf+5ydfo6BkNmLg+Pog5/w1KnuOKuMwTMb
lB6BU2Q68h+jRijb40QFntREZ3hctKVeeZKPx1a8YzaJajyXfY2P8lDBfF3HU6hl540SkVLydyCB
N5t8F61RSYAztgiOZbCoBy5Aj37+z0mw9xpq+WmrSfHO4in2o3hoTAlwdP/JNJyZAUJh3mbU1Z7U
DfdHRA1ziR40sqvECG9YbVlDH/2PG01b3Zc+9mXpWxVzJj2prRAdTxFw6S9S8T+QDShsw9DU0LEM
J68h2gWUoqhCBYfWCBq14Y9+eGyUIaSHwWj6Uf20CzVMSOlyxm9I19/OV1mBFXoKuZ2bBB4QO0PJ
RwqHoEkLNZPHbl17AUF6xrXLAf3RvCX5AGgJxCEs08Crdoyh7YIrVY0BfINA6g7ypFe4zz+JNmqa
qhzZhV5gH+5AV+8V5biARaePTqU6LfTzBUYfn3EqecIo0IXr6qzDgreCNI49yL77yCb99ExUVmWV
KRtCKHVdOziNTRsIJY7kOoM5OL+3gE7xLJ9h2tKprjtM18XqnR5Oz8ilLHitbhWrBO2nxZjWH7fQ
Kdlz360usp7/row91m4MVuFR8eR1SblLLK/Y4WQMMBqZ3NbfH6uLkd4gxMXUTcR+7YRvQnh9Erc4
P0ZU6KVKhE2RbS5QiKdQD7Srgwcd2s7FyKHQRHwreZ7Wb8MGssh0ndcD78DoTmPJNrxubuiXuaR7
pVdObK4UBv/3ChuVP0Kt+GkRO6ce1fIqAvlpo/7e6CiGL7vJi5C97EnJIikycUKMnTkDE0z9wHl9
lJhLUD5njdipv9BOzxLED4X6eL9VUCCugCuJKg5QZ8vWT4mZ5itG4PL3yeIP05JoNuMBuiv3hG2b
6pBqhy8gDckg1YqP4rOZGt/dyrmqXzSBAqtsb6E6ZpOIiNCmEdHeVeA8pweDnEU7KHOR9Tk8CXJr
gO4a4bGPCxF4gyQDjh6ypOC65ea2EE20xfppgzdAnuiGo1L+pvbGPjlq3wz1EN7hrFAEY/WsjrG4
DPZLqRLeMLsI4GS5fu1rLSwdLO20v07W8z9PgCy7LDTWlcZA1cb0fh+LVjV6NfWNOThZyiKm+inP
hEpeLevp2lq9GWER6vW6rN6UoTBS2bC3iaRLSbDvXjeVPNFIaFcoWjI1zGneWucVrEYjPL0soeQ9
TgMCEXerk4xT8UNw7IAwhpQKI9i474dmTMvfWon3btJAQGA5ixgoiI8r4N4xoHE9bLDgHHTAb4jo
MNW7Sk5UximJoqEtdBYvIsXqo8ZEX0frJlTIHPoPVzlZRd1/StL2rgWxK86GNRcCwSWotXPwF0AQ
t8COsO/R9JvTvTIXgZzkWK4OHDhO64iOGPvntIrLEfT4LsiIEdmcOnCDQrxTiFTDFyfJT5yWtWk0
zuc7mWnUVQ/gXElVTx/K09P/Z6Sa4pTa8WqBJ9kA5bEvQ3WvQQ+CdKIxR+ldz5benm3gUB3khz6T
Vi/1gkwjvNDT9STUyJHaP/QIPuIaNEPxzhBtVrE5+BkM45ScNoV+TA8ihXEg3Da4ddEOqySvIkg6
g2h4A5JSGd4+943rGh0LapldJjWdfrOttuVcfoOAX4vqBGEvvr9ACpCqRx0L40jQ5ucZ9B4QFrZi
7sTqovo5gLMQ3RCqcXG9/mtTh82VauMSrCM4NSNo+qHK0A6fw2jcir35B8QtNx5IATebZJX/JgaH
dEDhI9/DCIBbCGZrZpCeU/Jq812aY0I6TGrPGdul72zZXOJbf4QkuMONz6fmaEnFhYK4A0Q83bAJ
aef5LsaqybIzo1twJfbM/kAR6uMFEXkcA52ZW78tkLr6WQ+QNmnlTVbgUfvul/ce0LlggVKkBB/C
njzVDCMsSBSHfQdNPimcL4dCY+huBcqb8roo7CyBp01DsOfyW6KgZuYqoWXPVfQuXsAZ/HM6XR+r
HJolfixYn35sYhwfxpzVkZ84oo/3rbrWTEE6uQMMVNg25Wcg5Y34FOBQjQ9uijpM/gjDuZoRP3HR
HvO0kww50NvwhEN2Qk7hSvsQ9KxWk+/5jSJ1RZXvHR35NnzQMSiHV4swnMoLouuSxOo1Pix2ybj3
rgJ+7qdhDe9kL8GlWeX2Hyk1j0gZO0LQt7pckA5MKi89+6qBZ58gu2m7YlokHBSKGTj32eYj+DER
pxJWNJLfFaAh0t8fpZ1RKaSkLKEKiznT7pBpyCj3myXuI8ZV1QJCE6d/VDv0V/wW0NteUNyjlgPf
qWAONDR6DaFK/Rp+aunvJ0iAveCnTeZYUDdKn/WzfSsD6f/jqtNfpGwESym04eG5i8h4KY+zjF3F
asDPIU/0SZ4phLMQUaZytEAaIt0qh3jI4BEvINxxOQM8Hmwgo7SMAoylK9vHqMtyILzhMmRfx5JO
fuLztvXKHDLIibLyX0NywCdRKyzYrafkpSGPHDWn6Iz0wkocYCJqhvSR7nI0lloNQZL/jS5dZLHC
u1dNUCKRNjEDsxHgEiGnHVpuO3xx7+Rhhz9oD7l01ARpXr030wWm8AbtRa1jJ/QIj0r5V+GeX5ks
eEoFSpllKNDiPu/Vh2UAJ7KlmJTzUFpYkzdAOwrPt67P9NOjv2/7vpJ7RmSmw9tk3FDgxJaqPB+d
YuYmCpETg9pHhdS89JPhbIyLfWkTst68mhJB4ClwZx83TZrHre0xNV7hhJUVx+2pBFndEnxGuyAN
kZTrs467Sg8Zlc2Aw4St/gXj/afnw6W/AUANlygTWME1MpEmTW7zCv0zTvykJtK0bmKm63EjPiMT
ZKv71H58T3OAesk9RGfNfzNorhFZ8bR1PiSm8fbCShl+R8Hxm2ljBp6oqnK7M2yOqt5dllapg4rR
2i9/l3NAaoyn1ANF3V0DX4kuEsgEJtWAlKGMsCIWcXtSSW2x287qNvwXZzQX+DbA+LD7Ilz1ciWT
6LdevHRpMyjyUOBjzYuyEqHAdyBmkoUWdGLFtggHqHsB/fl2LfHdW9Wo1DisqH3Kxl0wIXyV/XwD
V7gHtkUYw73LLEYGXnzckWOBdLpUhrxDrlIv5Jxj1OIjpe74nTWDKCepvZ1e9Av7PhmXfNrmNOEP
35G6wB4Z8k3ApI1gMmASjACiI6WPo074sDachNWR7RcWS4nzQitzh4RmYNwv+JGHaQriL+pkHHoX
mHeS5QdJBzHBoVZvy5PZs3EHZSlZKYbFl8ta9/4vpKm/dycHXiC35NG7zFlLK15Ol0OzaCnSW8Aq
mOqh84zjmgSgVq4bnpb6zwXmRKA5JN+JqyAwsX9juGJfQszwqnaFfX3Zk2Hou2GLPbT3InzSjkD7
0VOVaXi0Ak/H/qKTj7gJI4CYCUu8snK+CwyRY15SWnDLsswwwp2xf9UVWTJMo4PI4aOoek31srO/
187Bbp4PKiDCucPIVjt9PgpCMf4X/4P1EunB8BzwwJa7xywkRuFMSUfE++8xm/3z9v/Y4uoz3l9z
qqOetcRxIrqE3YPYu+jG29CKqgDv1sMox0oT1vpWLvJeo1D8ed1ADKBXey7051kchnyXTsM7g35J
FkTpbDQ2kVX/1I4yRw+8CwPtpS0KEgzU9u2ezsrFiD7B8KO7+LECGa5MlS3hCWjnKGkVzrHil0v6
uu/1oiwOtTY8tQvf6/vo1uGVhKh4NFokF9+rEhaKy+DVsY2bD+UH1kFXbo4tHB1k7+0f4dokN/Ec
dy1sJPs/hOV8WJ9Z10eWAEyJJfH4JkxeEn5cJuSLlhlu11t6IBYOtcPgaBmMpTXfQukwQVEQcV5A
uYFFN5fr9bjKKRR2LUW+2Im4YD4VchyMKmLqNJRYh65LFtiGv1UOkCBaw2RhQyaxkBb9chk5nLa0
JB3m+NCW0gCC91Iae/syf5Wtu4rzLfBlpHdaetmmnNrH2VXB9E6DeJmEvPyE+QkQXu/QRK6tP+cu
48JFJbjzt3yG4uc+kTo96yIGZcCrOJIUjh4HmhxcgPTjCjzwO3/0nqwi+HCW84vK9lWw/cUZUVMR
w9lGct49hB8RuCgMhYxv2xx0NzSNYm/I5cruNvSapx/bV1VCwlD/AWgtYFaUgzeKfONyzvAh/vm5
RMe8pi+tmq0pAoWRigAPtgF52gaPIbORH6GNaJGe/2ZN+l8NduKvRB8tLmR32NgfSZm+Z0Le8rg2
HE9OLMknq3F5hh2M6C/qctHW9PSU3WfXT590q161uHf+DCmCiRiB51Sr8DBdEx6w3knkU5lTypZn
ZA+UjGQq4bz0fO8Wu7Wq9ZoQ3fu6exI0SGJnLqNa3gSmgKOpWupi+Q7CcR5HqAQyYCYI4Z4oVkhZ
amqIjhezLkvzCiOCePhtcNoRFrgv7OLXHR04wG5j4UmFoWOKg30YvPb/mu//5nUZ3FY3zKGf3SRS
zOaUO56EXlzalMTicJIZKcYKi7dX1fFdOBwrvc1eoR7r4ah+GJoy29ajpwOJaHVr/Mxc8bbovx0m
C2XIFZXTG5dcb9ymoWVvrqtvcllMbsA8aKXx9qBaZvEjQyox/+zmJ32dtiuW6imXw0xHF+dvPlsg
ZSRrfbYutUzJASEVdVq3S8nIpBhuZoESMT51gk3FgSa3jhJJWF1nyWYyk2+V/E2bfyK8XXBlpTIb
kFK4zsz/kP3dRc20kUQnfv0AbDT4tigLaUQ0rL2i6BqLuuCUIeBWN9Uu3oPgSjfNJLOgLg/Obhda
N9PSpKTpR+jQQDR5ynCGxE/SYVBI8bhQI0O76fXW+vcSkbdAaKebHmdzs7wV+gqKzDCScUWAdxbO
YITrC0v1aVR6aJ1Fv21N21LQbhtnRqPngIU2Z9Hd4/xgR7+TsGOp9+1bmnbteqh6Brl7qpsmEPuO
Bbld/r2yLRBDUtwfaKWhbQlZCKCXbmCIUC/lmP/8V1U7LxmrPBTa1k9YsaF5Z1A13ejFviIcm6tv
at1y9j/qJjE9yk9YEJNeX0BdzuMqtZA0q550EHJiQAi2ajGgRQ+SYKNFG7VFxnoqAGJZ1J/Z+pDD
SSw3nUQxFnXRI01U2QQn4p2MVrAdMD+usiHXc1W2+bOhoDFzNfAtn43N0nyFfO3ygLhRuHyNeWiS
0GkgGABbjqWUzkzKuPfhJp+9dIPH4ofKwpIf0xwEXaxAP/suW4No0Pnr7n4n8hCz0gEWivbNOSol
RPPAa9Y9eaWIyniV3X07qz9oF3EUaS010rLF1MgOAT83I4xStQgtHjgOA3WC5XZAnsCGypsU40ZR
SDDilc7f0Uo1M6t/gSvq09Szll04NJ8EL/ounG/H5/PdWpJYGNimR+I0M6NHPUXp9DigDY9tGCYJ
peQz6x6u9tmZ2KN10ieHqWtpBWjmYmYpmSOJbMsI/IwYcYgyY9e5TwOeeTuhohiOgl8CoBomCUNJ
5HlvAOtTgBTSdI8EmBaAZIByv6MZOJ4EVNQ0t7b8YN6ABBJmVOjWVJNEZkn9An/RQhhj/XLBTGNy
rtvPZt3TaPbLwNYpdYW1ULOTXo8LN9ntM+iS0nb7w9NOQFwIj0uixyrOvAxUqff7t/1kE92oOjB9
Fv7usGxwIIaWc1yauaU0x2gV57y0heU7mkcy5F9AY73tYBHer3xU9h2TURgw5iqoBAvsl6rj8QOg
e10Oeo6khFfohVEPp3Tha9xfWZPlx7RvylbWJApootHrhrXW4xUMM5aaS4lQwhIneW0dEJSLvhD8
8assTcNrzTG8o5rHGcGTHTC9oVnIuwcVytmdaztUf0PIHI944Yi5sBMxv5wjG+vAOWqzLOi+yzsM
OjdxnXR3MN4q9jh5ziZ3zuYa/s11g3J2eZc0nCQ9XDGmNMjKZ7q6Xzg4D0cMJcZfmhmw/jcbxzzR
AtBIvRX7yB/X/m4pq7s0uvEx4KwluTyJ41OzEc2LUSgTeMRVUZqtJTTBAsdhD4yX9hWyaFZWGb1N
R4ebR2FMDE6zYMCQ28581je+sL49K0Ir6I6wMvxIJReggznAp6qQwRdtsQkv+8Hv/SeId8UUeS1s
bkj3+FwbDqIO+ESPU4yJ3x0cdO2GEXOj26HRPeX7mZkF6LAD7nPf2S0ouu0Vyktlk+mftZpPKva8
fC0ZH8YXI+nPl0pFbPszsrAA0zVI5krsOQd/pfIjfDFbjxFwtpPdGtq6bZYXUTSypJgGNSUIn0IP
STvBpkIsfCm0i1ReUichWJbmnyAT7BVu6YgQULer+Ve7QoVj3w72LI7sQiPQ/TA9GEPyPEg92sD0
ByD5w3I7QZ7H5vDCvvWzdKrfTvmg6LG3XQ5OZxPbXSzPz+7ZtJ3l160GlqJoSUONDcWduG5MrS6z
IGsaR00aOVVZqj+96s12blGv9Bf14Kgc0UojgFqIxzDzCdfaYvhsJRFpCjHTWAPaO4ojeqMftACg
nXadsd2kT++EfHyJ+gebKVUdCcTULPopGMb9seBg9GcA1b0sZwShwvuH3sHmrTw6nZ5TozUDlCgg
MzqlPZexB2AMzeoJlrLYE9EQzQoUzySQbb4W3dPoiFuM2ti1iOcgJpP+Kngb46ZvguiSHQ9gi44m
T1DFEE71GTvUSg6KkoV6MO3kLCPq642VxV/GLP2kanJlkGoepwOBrprA5ZeOzUjiAcrG4dEIDP6V
ohQdpvOM4r9aMOiN8HhlJpxpYbK6hrBC1Xjl6YnEh8nYpYIp+YeRsE1vye6g6D6mVhHaQi5aLSyY
QPFTowSHMwRyl4ENHs28r533s2bKXz+7ax2FnmJs6h6cveajfv6l4INZRD6HAlJgL3pEOuHR6yQL
BPMAo+wD25OSBJ8hlnHjmXZWmQh6hPHvzrxpQenw18b0HefnpA198+6dKXFbM2yQv5dShDRb1exe
owPuhtQA5uHGhtSTAkf2UvcV5myHj9HUCCnnElJKRx6QzgOq5Al1JrKtuccJr8GFeBKcu9tTto06
eNob+QMxAPCeaR6tZMTAMTvy8Ht3Z1zv6c8r/mU//MJL7I0OgAPAkb+JwS3F2K7aFGmCBn1wLtAP
82Fc3Kk208P84uN0kzDYlxDTj1A5A9gSa3J2uFccdIaGeGNhaR8xxKeH4Na7jcou8gOG8+xqfSxY
7BRw1/UjdHHvQO9nR+mpqt0aMgLjRu8fJaTOEx9xz7SXmk9RUaNDQ5lPZs6/7soNjNbZsIJ1qOWj
IEARtP7TzcCGrAMD7j4QYwGZ1PbYro4Q1YfLHJdXcoFf7nl2QoacgFhxdP3HY2KRRJPsvfroYUrH
Q4xB1cYauOdkLU7cfvPHAJSI/Y7z4AzIeQKGee2d7tgQeJDgmB68pMiyVy4LUYfZqFdpUh3slI2d
BGTNwxCw1OIAoCz9wu5E29dQv53hM7IHVYyP2XE5aEiOlffnAw9GnZbXW/qs4icfcA6gHqSvpyjh
gay1UFgFQWKrw9c0Pxb+HW36r2iKdvNbABRu7WWsvmbGGPVkR00fViBqjtOdZeH85EbKIV95FHQT
5kZdyJVjiUh9f7Aa0Jb4lCBuZAoDl2garkreiHGNEVOHEEXf0HRXP/MAXzOpEhjBrFA2j/3c9hHR
41jnDFhzvA9m+Y8QFmS4zI7qNLK1IX48yEKRtLqRMjScDz4h9ZwFVhbpnWMfMEp8S73s3BhBjYmb
xM+EmKMnhkS5PCvPJF5HQ+TtqfIpX7ff4Vm5jWn8xDQj0QtCEhCPJj1oeDjjEYCRfD5DU8Aleuo1
DedIRgRYlzuk9c+hElMseRfnEPYvyFBucRSCOMwskQPc3JOxo87o5IyHc30mIlwII0ba4g2gMdf5
WTevVlK+tR8+ZQVyDE2+VbFtaLbV/KM7oQuz3TUokl9XjU81ojsqB+PlqnV4bbfcwHLRL1P9Gh7h
7x1sOK58IuU6B2n/HAn3LEboxuRDTNh/H84I7rxVxpXpjc7FOiFxrGAh6h8ir2A1+TFCIzmKV4NT
yr7IDr46ZQ0blvuFjQ2NvX8PvXLFJ8casInpiYjAA59tVjJUZCH5MpNeBosb2SPzjVWMP9utqrbQ
Ldn167suxqaNnMYgGGenAS02KPmA21XWgz0TCBqQGFxmehGi2fvfWgRfN4NJ7pIu2yPZhybIIsyk
yVAaeTYrqpSnlepJVdKFCy5vHAQBro0SQDkZ2Vf/e7qeLtAof90dZxkZ2Z6PXgNDSJbqwoaFUXIG
qjAEX8+KvD+Wc3vz4NKxoNwR86+LcM5ZVzjRN0CbV6exhyuRNm1b07U+WUWC+t2U7YiT0OtFGciE
bhOLDyGMXlUn3zWXh5xQDmDuzwFNMpEkfDiu0kzjdK8E6Iyix/TzJnHpHCsDhUnLG2Y7+bWIHHmi
sKcsk43ZLjQXyBtUmLV2bJ9y0kONKWZdlENBlz6dPXlPSepTY/sxcror5hTF3GO8O1y7BrnIoRck
Q857zA8aD0LRbDGdr94qWVnRyEA+zPjb0fnLwylJLUmoBZ6L3jh4OWtvW9nMBeQpGCTEhpQ2z8K+
hCqu5S95GGt7K4yozFQz+UuYOtj0ZabcL3eF8qkW3NjTICNOJneb2Z9noqMm6y7mQ5nrI3xYwsu1
RypkEM7f0THvvFQL9upkbiaiF5QmBfReyhcarU9uIYB9ZTWQr7UjBJBtwGKQ7yvXWL78MdkAKgNz
WC+e5KW4hN4j0GMGgp5cLMQHaQz+XcXZ/RDqGkbKlmiP+Snns5xqXnDnVBAfMGtiD/dyxXx9ixkA
gUM/YX59jTt//wz30oqD7elg7YwBjWWRLEJN3wb4JD9kA3mTVXYCrNLCSQuuddZJtRgSG75mk0Cz
HTg2wnr0OHG9M/8ozUzWfacGXyGX8GhnLCLiFAaMsj/uaRVuvGt57ECpH7jGLS/sFfRac0oXmCjO
FofygKq5gtaPjdjW6CP7d6E54vvLB11HuMGIzx6/flI5GlEDrlU3P1jNjnW5b+7N//zhSg/RQtr2
tFonefAAynZKDMea2LpN+d27N2nl+uFCG1OUfIdfIg2shie/2sYKv6EH1MO/1LZmbAG3+jfC4PSz
qnXruSbXCI9Gsu0qo87OXzRylN6r4hZs2pQNT2/jaJS2P5CqrtOc2oAHtSW+WrqoSAhrinVijlLM
AwJ/eH/jnAuoOdedj2r/u6UdaYCpwEnAwmAVKEFXMqMejJ9GhdZVyRrNBXZLZciJziuLFLMuj99W
k/DTJE1t5y5PMmlYZvBxMAntDjfe/8X5WaulQf3IG4A7jW4YiSz3gBKBrhxWliKWMiIoNkc8xG/C
LGnjbgJ3EBo1tjuesNnKIrerz76wIEJTNvHTsxtobsJlq8JOq9MTR4farKhePxFTPJauByQwK4NG
MQ/HdqDFHQsxPaBzdKo8ppO7/31pSOny0VPa77U66iOtJsbiuszljufCDo9pXRwrOIc75LffXkrq
SZkQf4y84F+kKn+NgpkjAnCiwNAbVrtsI0hPw41uOrxwEQnJ570R/fuU6QR4LgXhEuUyAlm4pnBg
Bi4lEHaSrdYlmJekLPFBmgj+Iv66du6ibJnCOssAagBVVAn0EAYrCcYWuhTBFv5qnPBL6X1FTGZL
jTgH8FN94I4eKd/WLMCZDZx6yp91xxr2dE5ypW4TcqAjQPeb0rgERkFcgodr/0mck6f9O9KhLWHN
/mRoLJCfGs2j+kb73LOnZt7SC8YQVOjPAT0QFOjYpph/1H7MvPGKlsKkBcbIUuLbkAYd3m1k/+bO
bvMgDygtINapO6x/aRNDMGdA77hkEMlc+GrhtueqrWpiB+NPejKLLy6oGKBmGsdkSN4+Xao7/Na/
aIJy03SUfyI4D8jHhEOuy3NBNxCHkKP7BnT0o9PiNYqSCUJV/tNlOxvF5MUBMhF5cQX2Hqj1UJgL
uMOGMaXyl7XAuNDdmjFd9eZd29pWO1vuNqvQpwzYxjLpnRcT2EvW+O7c3OMEaLJIG+CDY1qt1zG4
iuF/ZAc+Js4bCFr5ppWbzOV1xdbHzuhuRHbPJcoxam+S9E6dMyxBpQXyNMK3jGCiLzjoQwd+E4I/
Et0J/55XxVtDamQN+1hMvo+2nKTnHTjeonc7aoxI5XuXxiHjrxaevRWc4pQP589Z95kMldN4RR16
3Z9YGIKovqF5OobcPE+Z3dTrsqHxhRvseZoEawa/sH0UO52EjqYbMy0mSvqu1uUeA1+OhRmvAsD5
fjh80DK/dRa1M5qJLoZl9TgOjAgzNs3S2zE7OaS/A77LI1SzUi45bR9S31GU23zg2oxEZmAuxsRM
c3I1M/qczwqttesZwngasd/dDVxoKS+9KWJiLI7CwOFbuBm33nA0fIcDBvTb+s93u0O3iQ+vwUTw
HUomUlE4rtPEtbVH8cCt6Cv+m0rQ/HBzCgPjqT6ceoQ/UiKMU3cIMEYQNaCiX2VhZ3AOhrz9fqZf
IGH7zM7BGmnWo0tUlb+SoLQJv7kP1SsI7Yev9Qs1Ky1HAtd2aivxVHaCc+KQCP+sVL8HLaVe4qpf
P8PgtL1yBJjYYVLP3y/bfOhz+k/kLV6eQ1OGzh8PuSQG9pysyZXyfEac0O12NQxVDPwqd56wYuYP
EQK24MjCKTeLtAAUgx8sIlZ8TjGrI/qEixmJ3HkZ3obcyyelyvZkxep+FD3J0CV0o7hsAA2Uy4Mw
Dp6vcvaSJTzm3dYutgf1dsHYB6w+YkxbbtflgGTYH+Uo10teMoyIo7gK7B1VAVi4nuKpNi04ty59
LW939FJSJT6l+8kUv7lwmuJhETnOdjjcSiFpFrycRdiOvA/E8bwdAxfA2RAaZ8ijPeOkXwPW6AZQ
rDyiM13srjlpl0fzW9gFZWqp2hEAQAdlF0pmofnE68P6LsnAsfyssXmG+XEXjXjeY1lBbEB7MH4g
/soTKoREj13UCT2+jBbutW0IR0UqHJZjkGFOy2r2G8eDrJbdIxgv02MFy1GbpERFUCaKigl8bWeI
wZv/D1iUbLfpqZDp2i1/Nc9n4fHQgMGfCQ6V47cRiwrN/4OIMPY4hldlgsRK6sZxr65ZFs6albPK
CZ/aAUV6Rs7dKacFDJ4BiIjEdsmBKXd6Uw61mrYdRF4+IV0h/fME0UIvEz2vvMgRYIQ3exzKTHnm
xOMICFIfVISvAQ7xlKCDVns4lIVtell6lsWXGdW2AnHFLmTGTpKnHYgeX5TscnVL33sHUKxwRvIr
2wHxQE6nlmq7wqr4Shpt2sbw6Oikf7EjuAQPGgfekpYQ3McMs1TwJiXL4pIlcr0T7DGxgTdg7yVF
l/fFJbZVDUuUyP2W87Bei54/6Z4QCZ6OQDdQSYEVWgCeCNHssJ0ZxbpZlomDWzZc2yPWa7Tu51qC
hkPeAYUhRfu/jF5xwmKveZzTbdUCB6OpVpww3QWc+d2ZhrEa042zrJpUQozwjx6xdXfb/1wZj8TT
eSizlmmuKuKF7qBQwsjxmSHbbarFYjre+5r7kxRGXFU+nJKsGnOrmsnmEqwT2ETPQlFQz1zUzoV2
AxYWFdCAHn3bb5wdzaGcVxS4tiLwlRevOdenvMf6mXFUHj3Ah8r29Uihwmh0mI9HmBCxzubwqV6p
sJZmu96BRS7+AqY2JLPi1AwdQYeHuwj+1asi1Z0HTpuUiw0Sei9F0CgfbceUBg0Tp27ikQSFUvku
bE8DfyfSu3d5pJtAhivvo3vXyTcM3hhY9Avl/76+sqhzOOLkFZzWfsarjKn4vXaJN6HT9PoyJT/1
XMpLsDwIaSGRQALqsbtcMmXwafKqs+3AminMxEAdlFIcXQytQUShdCtUDspci2+SHks2sg/HAIXq
7YjOPENpgJ1iEMmlypMsboeLQBTi3U8agW71ktDfGy6DE0bigCdhjqb06B7CO0V5w3AVVoCAL/Sn
HLqAiXs62W8C+kdU9bNNdQANM38R841LNaSYK6ntj9OyTd4GC4MNGhb3xtXfVqUrv9henVW+3rP+
ryYSS6uBIRTXKQC5zodzNMNWaYlM/MY8uIyjKlC+8kebsKwBXM4jCsVwp38woWqJoQEZARUm6jg/
K2MVI4015/09cTL1bKv/BMtOcaMUc+VO/4n7tIMW8X8sakgen3clp4ge5FLcvYKmf/IS25Hif91B
EoS740ZDkWq93adXQR30/P10wtv+oQFitk4xkHsoeDMlaWwyDBYk0VTdYL8JC4i4Mh/yZVdzOUrT
LPru9K2+inXF/FPgZwCqOuOtcgL7n4jacOnEYrUfuvuBdaXe591NA3RdaeTc3dHWZRFRPnCD8yKX
93fCrOrDbXOKCxVdZDshc6BxR9PPIE59JQFS2o0ttQ6jBB7O2bDjXsvGMk3m+YjXFQB6JVg+fD/B
KPjUy9rWEw0heOtgXDBy3vu+7mJmSHJlBhvdRvyuXL0zhDZU3F4j789deAn/37YhaBdvAaQ4AWbf
30WOCYJ8dcHS3gObyJuBhnUXlpHkCTYiqgnggPudBM6koUI5SYCKqLAGPFE9z3kYTEQYQeXYcYrv
7L+Q9Ic2ByXGTF+9rg20dFFIl3Ld9IOWP9Qupo3poO6ZJzn2itE4rZ4SCDOQD2H95NLpTb9XCliF
GPtvgLAo5PiSpetur4ANlLl7DT9TOJE/JSbP6MqDJRvljgNLgBL8wjVjPxldk8KqWh3vJ3hzm3kx
MdzHxv5sC7UWKT6igtCOfIrS8zp7iWSFIQ2DylvbxNFZxZrEjp6R0O37oTdwLFJz5UfhGOmU5CFv
HkeIETrz88/dIYVy9aUPCIvL2hR7MRJsd/loMqdyCQjrs3xEC0yRhUUMEvau9eoFL9lVRu4jLAjs
NcQ/DAHFkHHPxc0dMOZVEK44oSJJyoJh+hHJRba9XeWcyVEVx5wZ65CNAC09epZJRzgMaWjDVf+P
I9f+db/+MWqJ/hEomXOt+ET24CpneQUbm/VExFoa8bCV6HwC3V2M6P8dx4usMSKbhq19zA4oqcO1
Gq8a6EgfXNmR37FHT2LBbAa42xw7XpTgTKIvi8m6X7tbxmgiotkEM0QDV+pYsbOu4JBlTCCP/n36
gL+AfHakuzpJJZnECjzUMs0ohEZOM/KQAtXXBGXh9ZUG8gDOMhJ+asaVNSFoKsacauUlBgE9RbCY
0K0XvF3I+ApXlFeFFBL4yZuzJtgekpZCnKUh1K8vBdtx9YVpmkVUX2/qYh8gZEwRqERigZUCTAHR
mpzcEFNSg2jXlcwHCoyuv3n/FlCKb2IWhLYnHbRb31ksntXjIE9rrJtqhvnIKY9s9I1nbKAX5yg4
eJq545opUYz4iGEosu9/fz1ajl6iJx3HMbvO1rkjNnKonTQsbeWMAj01CEL1MPAadXt25clwkxN0
XuSSG5GtqTIL7KI9ErWtNzd8BxrUmZIBnj4visyA10nW+TvdwCAjZDW84mcKuOAmZ4RGb++TQ2et
UwZI+pWlls7iD/MZrZ1/08fZ3wulvblWdS4le77rBoLYRjzROmklECaV1SCkTXjVTme3WvIKrNZs
xwyM8Ij8j4cayW+83yVGBWMowpWe1eRW9oFIPA+H5hdOgqYo++WaM4OyI4/3rUCpgBgw1SJLsI5e
Oc+RqWBFH+QgqT1tWBWHTeLYCxGEVZP9DyJFciGeGJg0qOkjB07sHNWzH9kOx04kItahJxYWzBgB
8kg27xVnloRIE0Iv1oG0kNcHSUTP45OBXNtnORZkaAwbylB3nR2L24FjlXXch+1nEGBQUdjYyFGd
xnqxvAeOagxoBd/gPOhjRBKlXzBAheb2VfNXsu3Wk0ooqt5PGzKa675ymTzZlLPCEjOIS81ZRnPm
BvMUOHXnlLhW05LaC14UXZ9LUIZPI3pBi1iBJG5tBBCY1nAg/HmEl5OLRoaCG0oqvaV7fOV1YN31
/WU8tY9HYPTX4iXRATj4OoXubL8y7/F2HOj4qgGWocBAAMKFTkl2Y74NfStpSWpPxCdwJ2YFYWPy
AmiiG0zm4dv7+659pWAHseQDmLFUgp9iYz74xDzHisAvFZn0/jGTGUQW//EjgxP4OZGloHwIlKUm
OCPKhySsIDFEG4jiFMuHpfGuWGRHsxXLf7zituJdy2WktmI85U8/ycH/uDLVldJrPNxGY3zenYum
WsDtJ9iHgCmhTS9dYK3HFRRgWpurn4xEdWeHbIYZcl8z0cmEFr7CN3y+12klsufhP7bGIbTyDOaO
A6NBMCOegTQB895lLsvcLUjJHziFd5I3TWTIuWQIwa3Avt6f+8+8njHsaP8qS1XfGghaLy4ifFUb
MP5jf2VTErAelzR102pcvKxbW59ZESrhNj15V0SG06TQq82e9KrjTTr3G4b2zD4lnxAL+SxVeUzP
Ng/VEvFhwown/VSobnHp2eC3F5SsPl4viK6ks8Ln87Zq4+e2mz675io5/9i+pZigX2J+93D9J4E/
MavYYqIsaqWU4wgHf5zvGJpLaApai5ORzuCUl1ru+cYdOIgxlyBr0MPKRdeMTaizr5Cs7ZE4D89Y
Ncw5uGh7XWtjSwSqa4D36jStRSWKXJ579xnPnS3JYxWDp+a8GufozaJc9KhIecTvzUnIgHXitEXF
M4hUFLIlazZlGOJwzH4hBJ2EWupjsqIbcxbYmyC9wboa7yPR2k1SiRAdUKarIiOwfD6ano6zwtTE
6TMVfAfFuIj8RmDCieggAzCIrKeN+N/YhAjy5kVqV6V3aEnQGi4QOuTatvUzJ7pvF7P0qX/udEn8
qBv/1WZ47oxRxC1rej0c9xiXdkvL8HAEI8ZrasK8R5AaZUzGi2ZUpFBtL++vyHX7YOJCVo7bhd+O
9mLXXeij90mUV+XgvJswkZovNd0Ox3Pv8v4+b8uODCtyG6UxDJf/dRfZYucTwCmasCYhleXXo8bI
XgXUSslaAQg0OOUDKdgSo7wjcjxt/wFO2RKNjiRaZa0vTsSipzSpshunHbeXJ19YaLBrBjBPI0Mf
ulia+9JGROPDXgj7O3O8h95AbX/KqGfeYZ9JtwCCyW+HgVrOV0ah4N0jsXn+quvrrR0On+jWhD+a
aLEcRkzPrDaK7zL0/DPNfw2pKsk7+97Z8JX9mDH+3ivMV1CIaXxn3kG7NuFDFagqX5bySj7BK0sC
6kPjnvlmrjXMP8wGPW0qnMOwbnt/tRkr3OFBBquX3ryFTG/EFBR22XgtcGphEQuGd6bzn5IpD2Zd
TrHn6KZEJaUyXkhwD9ojvKY9eCAzgCJxXGuhK6RRa2Gb9vKvk1Z6c0+VeppDr+sirKI0HtGpUw3D
G0ZTSNm5C9Xw1eop7mDzCz7AIF7ZwlCVyvyFjUHbiU75NkMpf71RBdmdVoPThDCysRgep0e0gJDk
ZDKtRvXcadAOAO+LpCPBgERT/wk2g56rIvzRFU8Ca+2VLtpeDQXQWmI9qJGBW6DuJt9DkKvzd1NE
1yZwyn5zdf7uCVX0F1/J+AYFMdJrqh8hSi+DaLZYlS046vYS2DkY70ZQhSpEWi80pl4J/wybz4EL
LnD0yMiaEafG7gBQ7un3XIEUrext9UqrrRlGb69Na7i0Y+fH+0gH5dMHNHf5sE52j1IzjVcDbtBa
DdLVJMpJ/+g6Mhe5dDblC46hn/7KYNHSnkNQPV9JABhw3PZ8Aw1pHTyO8HRDwOQXyCak2fRBh6u8
kuATcm1ATzXeV2y9pQgBnfObwitNQnlcdgknypfiEHstQYrA8+GiVlWVsdsfCxyaMuu4DeDLSN+9
+T0SHfmNmn+0JC1/mUqrMhGZ+5tunEUBYNaaCdqDoxWK6CvMiEX28mKkZrabkETvuGKQ/2UmBiOs
L/dMioi9GxjiBYOCE6mvq7DiojCw9/Q1uSFA3yYRjCEPve3QhF8Na5qe1rBPJUQHlvZevyM36bNI
MHfoCjtTnn9gjjzkE/4SfDb0QlQxhYsaHLfxEarRid9x94mU/U8F1Mv4/2XK5xq8ekXi6At5YN6v
PRf2Bn8kYHdKfg6oKlH9vT9SWG1pX7HgNBxHHdgIUYAlSXLM5at0IN20Bz+gQWPrA/tW2Q7rJwpg
97q3qtzuA+p4Ar8Nqw9/AEA4VWEHYmpdpGFWGXbcR+DCMCw2jtACzE8HnIui8w6xYmfUxIQ3+bts
mCESwPdjqZJxPXm/ixjNY/ExEGbUD0xpMQ5246h3kqsipgJQr0zFhyXWLc4BelIIDEhSXZBgVo+T
xbBLBdLnLJHl7kcFqu8y9/pSSyUH+LvgkAibuFzrgWzXyNvg7Y2SjT50cl/eRIxgzm4EfJCJ1xOs
f17PoRJ4rLaWzivAaE9k+9++pCNd4sfR6Y7xW72QziVa57C7MajZO0rUftaz7HFPr4YXlrMaQ7Yx
Xm4Y8o5uyybXW8LP56p2UTi5YeDxYXdtcsu9chLIwgvIKRXAWGL/SzyZ35125KQTFOm/Jmy8UYWH
s0EXIebuFUoAJNpS/14A7q7Mc+xLrl6ak5V7ObAW4tUEMsYbD4SeN0iGuEVAEwENQUZ/b05iCJs7
eNdHPVKpshf8W8Wd08gQp4qGmSBLnREj1yZgfknyAzvz40Uqlxh8TChESd6bvHxRjChJgic+c1FJ
JJoI55YjUnx6Kqbr2JlP3V2t6oYPWJ+Y09cu7GPerqf2CA1QcqhWdwD5LkXXsIORxRozCtpLh3Sv
IPRobhUORstZdWznj02JB225AVgaRVpPCQHwvzwa6zwtdw8qSY6bF5xpMOpCHvniRw5K9HrmWVA+
lKhWRFXFMSw/7eWuc4IXLgaBZ7PX4zBPlq3IpbVQsl86ZbVnJcp8/L5o67JJ79Z3GHbip1AM786d
iW4m+pkgfoCu9rrUCE3umQrtWt+BcCR0hcXWRu9YfO8uAxrYdzwSBRLyWo77yy7b5XK9fC2xQzhC
8CNJk/cRMoxLi9u6QafnQSir9290wC/tUC707b+sGBlls8GkbssoP1gJBCDGxv2XZqsbvvqm4Jma
N1cRibqxijzCPKpd5gP9SFgZaWCz1hNr8v1YA/RWCPUt7F+aiUKSIq+weiPbSvyXJeeXv2ZLvaLu
dn6TnyDnDEvzMWmhLZQ7yQZgkXWG/jMeJBSSW/OIlB5U9Y+xSXc9L35yWH5gVXE0F4fPL7yYR45e
G167LZNg4KNSKZXOWXFbo6/UkwNjB4RbEIIRSts5sWK0+WpcdISiktUXQsz0JVhj00WS7sMMiJaW
W2LW5cSCeFmq0f822PG9VC82n5MI3y8kVsos4buKiWEk3wggvb0r3+iLccFoP0DkGNPizhRCsCu9
+z6AA5dPHLDAtkY1nZbsO+4L5CRkmfc8S8fzQO07zk7noJd/3vvJQoYjuT7IVDFdCBGzVQey+Dxc
MtTGAtoJWRWtLe2fL9mXq8LR9/cK9aWn6NEKvDcHcZQcnqT2bdQe5ycyt6QkF1dzGmxJqsCx8/OK
9VcC/0e+oB9u860+gtum12BM+3u2B+42tBE/pRAda1zg/QIS40mwvdkMYcDWKHJ3AyOb3HxQ5E/8
NH3xgqUsG2rN2LuXun8gQxzIJPcse9KeQVodnYTJX267aOgcEM2gQJi6/ZsRc4SBY/dCkl1p1Otu
imNXiT+sUBJ7In03ja9h7P4iZX7JhEkef2Qt5QX/OCYWm+nT9PVEMGZtU9PyeB/bcLq7G1LNwXo9
//K15ydmJWQAcxRSLDbJLxyVgWVmvJNDYHPWJjA2k3AydU6o3vbzMZFl0IaAi1/7AOnzr/uzg7+x
pRzMU0VEYw2OgJ6L/HLrmskV8o0fLONJ0BRvP/lm4lt70h0PnuNszTIYq8/CTTWjWo4wAiNOpVaQ
q/TyMNha+vnj5p5IwW16pXfkS5AKVbGqnkbb0foGpqRm14dGTr1nZailK0AmV9Jra9LinbyE6TTf
63Gx/UnktgD+EZ3/r9awNwyX02O2DeTLZNuK7/K/w+dlDqgm3mEnR7V6lawuCo15UFMOmPfMvRxc
nP3WMJKZGSHds5DDDvR/5SEspmW2iLt3BwN1pMqGMwen2mjqT6vekEfQQCAyB7zT/nmLLPbh/vKm
aJOCwXLLtWYJ4aKaWIEZ87871df/hl9klDraQcdT+lHmMR9MKUItD/gi8kxCp64Q5Cr6U5Xrwn19
CgYyF/OdaKGHqjxAlGwN9TcvrxbIJep3MAgCE+R6BmI/1Sh0JWyFjFMrIhOHB+0WUFU4gDfFqqvr
/nzW3nmYvCKPdu9m/S3gFjNCHQBPAYGrmbdcBubdLfWidces4TrIeXhWwAYl8YYTaMYR1CHjSpuA
kGLkTQFYbV063j1rLXe5CbxEGSU0ZenDDhXc9AuwPiYTBd45a8IYaEHZr1KJ6AvpurqyLS2CAyQ2
/hc7PdvwksMrreY3s/U0c/CyOam0cN3Jw0vRft3onWF786YIySfrf2HZgDY+Q/GzgUCG09PHw7Cl
L/8YQVOYiT5+BaaN86gd6hP72ENCFG2C4WXy5pannrakjNurlvONfxEooRBp53j0pJkjeAKIOvjF
0ztA3AJMBPqLWc7JpGsczTXa3vIawCbS4bVlKoF4jNazjdAR75AAJppsCJfoohar0OZeGJMKUoZL
p6ZK8OHM3YyHXH1gerpZQkG2YyfBus0n7f0dUN749CDgZcYTHJSDJKf4jadnEEUaWotdrAtUDcvd
QjGasdOQxbby68hll+HuKQ8ePAZNK0o3H04D9fE7Lb4EntZ3ICcm+AhmxqC18pFe6ns1drOt/Siy
kJ0ZISDyNcAGlWnPIvyp99JsN9nZT7+H8b5ka1GY59QRMEp4TBGxw2vfxaudbhPHpOvHifGEzfOd
qD3EYIBQOvzOs+eH8myXC0UidPv5CUIqfUY1KIM1hOkZZFS6LxYmjnEiulqmiVm69tbMog1+08LU
ozwK69jrQ9oYao5HJcLF4WbYKz9CeItUnZRYtxIQj3jjxWeU/uycqVzRZR116MB3wS3RV157E9em
+RXwT9so1xGgbH7Yv/92j/rfeCYQRJZh3GmMiiaEt+xu0gvYWN/aUPqBRruQJfNl0rLKw1If9oWi
Yb/VPgu7Oz1Fyh7FyNBt2xskiwlfn7833KzGRX7c7FOfQ1Cd72tyajuPUSdF0hPDdwuYDcTB1gAW
kLi/8rDn+ieLYwCWFbWiMQaAeGZ3/YooFL/XiHmjjlSE7xAdvDKFMF2RmdwdoAcIRpMCI2YOAiYe
kP69tgvnFUxVG4LochEorm8+FLn/RZ2xCTBbA8zMx/BzJ7HkMTWdKiSQ1CFLy26s9Xb5efZ0A66s
va+I1rE8Soh5SA4tkzFt4wVcHrYeCh00CjMOZfVafqDMgukx1Wkli5O6IANpYjne+wwycXsgX8yE
pM8SDyfwO8hYedSvxZuFHwT6Ehj4qvFE2nkVMgT2DtAtzcFn/3wnIFiT0eqz9lSTcE8In2f8PWQ5
g5xUxi3a396B8nO8H20YErgHXdOYIxoJrbTiiD11Zz4QRQkUpbVLszuOYKJD1Ks/PNF/t7aFh/58
diwbLPwEouIUECf1HL4ME0Bx+HA/Uhd/ukhlx6ixq5KDB9qzu8JGg5x+sYKKZVCwx3Vf2hlbp78F
wMGNiQrgpT4TbK2+HNMOUaCAQFhktTPyWJ5R8z6/JVwl2iyITf/NGdCimyA9PJiYAlPljUlvcmo6
3hoA3r8HzWDp51Kry/VmxB1xa0eKhsn9wejpsPfunpmOt7XGbXui8A4n/aa/jFyTbMN73hiEBLIn
SdM6JwiBjHLfdhX2qzwGKwQXASa9BOb4drd/zd7uuF+vGDqoMYCZDDkqlZmM2AB2301dzFcV6jWU
MqLdbUkuKSjAqXBsoW8Ct10S6GzRdVK8dkcePg9wqaM2g06Pv2PM4oQdnBadfcyiKzViBYhxiU4R
idDV7A7bwTorLGIxJ5TcSMGfRFzy0Ywoe9vwu9gKKcCQrHEC3XEmmTw0XkB2z6OZUtc7sVgOWAWr
J7aoSDWOtxdmcRFdI+AcOnTXbpETJ4qNlBjOT+tmia2l9LbaB9Au8RgfeJC55aKkpMmbTJS+J9GO
Gc0Cfw8okT8XaygNkC9v9j9z2yXSJPdDd+vNgXB25/MpF/xYN6BFisy18X8Qk4NA1R64ZKtJBTwq
4jdlTrr5xas15NJFUPbWFxcgmySgfkupfoSVef5z0kyXgVsfCAh5tovaJerzDO6pthgCB7d3qtVo
mOkzt3+xbB9zEz5s0p6CgVOWyGPvSRPRSRa/Wm6MVl6JBqCerfwn/Wsm9npoDFXGnEhNPFQgy9aN
sicsR4hcLJFCk4KtDC20KvZYsPgKeJM5SgwDp+wBvELMUe9mxcGK9puB9NDioI2bDxmzkiE+doYW
rCL5mikbDzkoURUiznsFPBw61AuJpGAv3AnvI/OJxudkGLksIwl16n6FX8pDYBFz+D+HwIlovWg9
9XoSIKxCMDnJJYHFYAbTos/1CliqKCq4lsMHziey/Xnzyt8YPTxrzUkrf86fNkfsPAq15waMOiWi
utDAw5n6gaCZZoAEmYJO5hBgslTV6yH1EQAuAfWUTMmvNDVCgz8w9hK7cNP1i0IrI2JLdn8au5Mq
OriuLiPJdfhlcW+cRKvuI5+C9KZ0ZVhO5VZt10IQPnF412qAaaU7rqAQOZrZH42mP9XmBy8D8Hj2
MC3f5W3Gw6K8h7hw9Td3T4hspLOuT3ZCp1ZUGShauQYCTQBBhnvRtQe6/CCuf+QqEDDIpitbnXl2
Vwt4bYM9Parg/LIDhJOY0hqUieHWvXsm/97OVUB/7uYR9tiCACrYl+14GGlN2RsbAX1tXI8j7MZ0
Q+OovH6LQHt8YLLw5Eew8hc/vX6H9REXDyjO+fSM0IWyWhAEAgr6vl6iiex0HDT+sknDW5cfo+aR
EPvCJjZUrNQW2uIzkZUhB8yNGPjrDD6X+id0Ru3+FOMQZiRbUGsjE5O6bfq+7EC7sobgMk7LvZkS
EbGI//5Yw7xKEUKXEBsDfOhPHimZt1H8xQvaJrK9oZ8xXhHnDFFfTdjRY5DlmUf9h9rKBnkRlgGJ
epdD4+Ld4oMZ9S82nSHA/TgYw0cHs1nRQ01136MAhXugWyK6Gt8YYBeChpPYNApygyW51YP7FIDQ
AwowihKrEoU42lxI/jnpGW9yl+Zkm6mg+42NUoY2RVCrjcCBaVDScBl2M07eQEsIZ0lwKgGIQ79r
6B4KN8zgDo/0pvA8bz5+resGP5WnmMmWkwgtUVHr66GZJPKgi60QFprUp+ozpt/AvHIDmAb3GkuW
H2KtT5F4CvPuhi6jLljYPnQXHIclrIcYvdcxK+YiUQooUYZtv6l/INqiBH9QlMqK4ZUwH2zx7Bc8
uyttWvXpGr1vTbaRphZMeWWLaQG9eX5YTidmMMGkS4fQly97XsZrTFTtbPja4+y518GSedRRw8gk
RgGs16xHzfk/G5MlLwPMtBRnH7ov5hbGwmWAMM+BrWsGWJRN1WYCKJRFgSO8aJwaIt9EMM94JEZk
1+HL7giiAgJnABtv8SCI62wktcvxRFTrXQrxI1caMmkhfrcr1HekKBhZVR5Mv11mwm4wscjhXUJD
Lxr3H/1OhjFCtQQE4DkmGZqPD4Jlh7Vp/lYwg4OJdbrp4Kcx5eX4ASFi4V58aP1ZjmMKU9r2FTxk
RxuKfHVcSdp4dt/50spLU/+Q8Ql3J1uBNOlrLSWOxkAx8QYcN57xRC4hO22xw+AJkwsQZUK9ILMy
L5mgYwpyYolTTBhcK/Tz6kyt3/EGwQshLjqQc6tlFNi4IKuLdZUWj92vvMFKqNKGDZSifJdD7PuQ
Y9HRF9LJxbDwnKdqOB2oDBuLjXiajvIEHzfjSr1J6jFulNXg5kJnT8t/NeEX1kjqIyBgcE8jthY/
ynPPw9lqy6pxdiYOeGRLu4Ys0w7vFK2tL0zc3AxY00oDJlqOUSETYgDEBeot3NYfvA928GEHK9xx
TQuSYo0MwN1K8G06TrhFVWKiPiTHkY+JeQxKdWGhzsBrYbO5WyebWVFxoySbrj2cnBy4IlbGGY/s
Esoy4XqS1Xx99mjPXC6zbyr2VJWGytJ3biVgnWgOd/0esG0cezwZttgUkwxvJqugssASF2tyNuqJ
nTlV82rmEBd4ElTrw7k1eC6YkKOGhFQHKUxFLX2icKXt/FPyHbSRPqdTp8yf/gMz+ooLREtAftXo
XyXHL/dgIo1FbmrtyKIFS1VBzXuhx1dZ1IlxOivtsOwMb7JbPaCQAvGianSUoamdV1x4g5csUc1L
IZfmSZ5B8NiHlB1j8lmBjm7F7r4fP4/4QVZ2me7AkvPgThmALBZzajPT0AvdfSNWiRAAQCKP6JKt
OIkBRK6kcCMeGQy3mvubCIiM3VUknJitjLH9MstzFenxf6LI3EG2BFswI2x8lQsRUclM7rq5DfrP
aQmjkf1qIHZVRu8avjgErRb4N6VGO4Npi67zSfGGoK2yPuzzZGTdpdmqlCaeQQK662XBpmgz530D
rn0sqWaST0ZB3syeS6/l1OjMj7ZwO+tI2tMsxnu3He4aQZpAxUOYTvGMOGNpy5G/btlzAMBHVUTd
vK2AiT9EuJDjFTUzacTVu2rNZZFUDCklRCDs2WKVNgj1MNAqWrQypFB0GcWDhxcuRnNNi05Eps2d
rwuzchuKUit+vrTTC1pedJYjpwyzi5Pvof8Vh4YLOuLuir/ikzitHsAw7YQXXrbjrtj4L5NDRgHC
GMZTRcuimPJ0CdpkZ06XKiyGizXqcshkQCDTGveNFHwqslec7VrmUIj51Zq0rNE4I8VvPn1rMSVj
VQMCs9vWupmLhH2j/B9ERWBsmnp9CYHcD8wG0G/2wKLuMBCSoq2gDAIcv+argb1R8hRJ+xaMnnWW
FDctLGdJwqrFUjfEe8Sf6uYHUkavqYn3IeEJpGj2kUJkdFAx2Vk7izpzLBZf0C2vtm9bJjPQk6ph
gAAmhwMngR2gU6ZhFh9t+BhHIjSRuhBM5nTDNQyV5NzDm4kQfL4omuZBYkMFcu5jNM6iau8b0J8w
Yluy5TJ4XvIIYoFCO6haAjprX0T690WdSVo/Ge/KqZGxbNofgtQyBtz+0XtCCLYl0K0U9l0SrGgg
sfeO2OramQqIJA7QEyI0bnHhw5kykz+1MIhDa9pIHWGKHrJjCGDIg1+o+0uECcUrsvE0PZL4x4YZ
k6u/UJWjDlX1Nzbp8mL7ZYRRAjYZAe2unjHPeuGvNP80qL6mR4vuyL4h0SuzEO+DKqr/+TLtT6La
r7k7cyn0Fu4GdzWdRo8XSmhuccKXsBiREbE8wTGqw9xtWPvZaFRRiFhxMKzgQCcNWsOR1sXMy0ZM
0YewmTkS4u8sS3WvOiuKHl3h9HvQ3xJ6ahSCwCessaUEKjOAZGCfYRqwjF1Jq8JuUihS5nqr56Kc
grxYUHACO4VldGpkpBQf4dWVJniwpz2uQCmB2H6KNGNjbtbt2GatwFoBzY1dOKkmocNAJCmBTiQd
jidxRnTWRtswKUfbnwJZCCJlKTWHmobxJqfi5+pntKRJZ1J14aTxrvcqzR6IP2MLGctwb9OYrS73
ypEYhAcD20jQkmi7ofVCtjt8tz4Win2xeYwKuNpGK5zDljO2gImPPzzQ6OW+zsG1nmVGOmLjVl6X
rVC7cdgGGcSZJmi5WkPd+QwKEX+jxmBThF6PVWXTF/bLHPEIqCt7dlUBNSCF2ehtTodwp/8YJxII
Z4EX0wEKdOUW/8WosTf7NWO88wU8S1UzqLXTbmtSNEqk4fw/SLH3SxpikwHh2V5SNSt0zY4aBNFS
FuuUlLq+gc/ppSieXg9V0qvI6WPa30k9apQUGLxawZA9VBmm3ILpKiPbgEIV+DiUEbCpG1QSX2w9
gPnrMgSqX45XM0pwgQ+0Dm7gITB5+aPTnaX9U5fs+kcFNvQQn4MBd2YWEs5qFWXGkRC+Ts5kmk3h
VOKXm4OKAJ8983zUaEpgtOM2Vqs4aXZnIihrocx5sF9mofDkP+JqbmQpZUg5rjNZB8TIaZ+Ce+ny
dhxX01M8WI0Xbuw3EtvVEtXFDgLEnxU+voF/PQe4FyKhVa62IGfigtsolObbCuNMZwUaRmLS2T+0
VBAvjdovMYmhgWb4QN5V8s3/bOq+DiA+sDeSZeo7Qkj60EphqcxVmkPDKrfo6Nu0HsnISALAjhk9
kRZbf/tDCo3j+6SIXWORMWBwuRS6ctcbNmbX6KH/WTdGMFQnIgy+aWmf2s1j47KkmFoEZIozKm+t
StTRmA1ANEnNq9fqLUABAIM8Ow045W7qJVmA2aL+AQ5Ye9BK3yl1Q03ye0E/gg5XCi+lSC0xny8I
MSGBrW1BwyQ1rWvEO39fVhQ4WTmcQwWnGLP0yZR4FKAO2xb7OHoezRm821s3VniuRVTdedTKV4Bx
MF3LYG5hi5IHGl63eWDNFcbkG4MQXYwb4XfzrcmKtjkxANLSDB0CObgM2Ln77fRgfVVc/2U5YTuL
1oeCmE7hejTRn4HHL2AB3E66dIElJhR5KomU1E0zznYcTxzJUqJDCRe9qHAcmBd7wxfIWugCtDGI
wsogoegypjYl7ujTYMm+GOoR7iototGChHWHFw2ju1Q7MqUtE6PbOY5FnFmy20OlfCHkg3tAyjlj
tuESwMKUz/VnTiFTFlcu0qGt2Jv84zuzFBCfK4jMYEIX0W+Vrdl5Bq6dOg0KtJOqXumJ27t4Xs4M
+WZPV/WQZmiZ0VijeCoevGE9U5GP8OsGVX2959K7sis5RLND5yYC8zzyYs2EmJeVljbVSBAB0UqW
2XM/3ibDeBD1Lm4zSo/Yf6AdghZbGPKuZqkiYdTzCja09vOXGbXJNnHJ0o/UOVbnea0kJIpdjxvO
a6jSvYisHw2wRnjW1gDo6JcgCZJDUK7ZOECXCbDUfUX6MulX1MTPb8RYA9dlcVwDeW+w2rq78xJ0
ee/OFDo9/IsxLiVtA8Tj2g5AWbIfW8H+g/1DVM8D+OSou1gv+miovDBieVIvEM6FpuZpVdV4oKz+
QynqYdiGXrt2jLgVSWQerS02qqA1H/Q2H8OIKZBaEYK2ETO3/J74V7OkHgqQDN5FuVzyw5leJDpX
FVnOHtqiqQj6Uns01sR3BYeFdoDRPz8eIahPRlwYWxlw8n9v6DgHuW0n8Ff+9LEzSKtW1U8KvCBk
JqJ0lMbBqGh70LBfX1dWAhFvM+fammWrJ8DInHok1lvpOPH/q2GtAGx+8L5F1F1T97iPhShY8ICg
2MRts8kWqMzGM44rUnHRXHHt3uAR4P0fYnE6aXftC3BOuGSZVorBlpkSIdMmztH0sYsdRLbZUNMB
/UFwU+oq/5YodxJ7kctKiUPrt06dAf38qw53SH7J5uf2zWecX15F1eIriNhhKAvNbAAiPo/MlZim
cxZFH+x1f1Ry0f0RSvioBEuDTzlSiMK73Hr9y2Km0rF1v7vad//lK+6ceWbvmfywegAP0GGIod0A
BCv3tZQCaVYJITvQA2DVUx+mJfvpR8/04i9sYyXdg5zIVoAOPTAw8ybeE+IPXU1uTnZ/Enghy+ef
gJAYHNeYekdxlx345vT4ZP30q82BJw7glvVZto+gIyk7fPxAXOA+EtKDAN747nLohLyOo9ccXCtc
aw3r1g8GN1oO7t2JkJo7i6P60E7gd6LQ30XC3dBMb0csVRQBoPk/S/1apprHByYBa9qs1iGw8bkl
ojeWxK1uIDloJBbP5qI74Pv31lLyuytiLgN+y/EKAlwlev8SKfY8JBx1bHjrTfL9NTBo/VpWmOad
edNai+Ir1xied+0xM/pt58j6xl+A/43IM0Acz89zvmzh6XM9T+1ckiNri2mDTgF48zbfKJlKDyk+
3Yr6mZiEl3d346lWlWkIEKvYKXeJECeqlqV+YGiThFp++TWNX8U9Wb4ZgW0b7rlJ5od9gBMwXYen
wMH4Cs0QKHXAV+Ab4Axy0EbdNvj8A3+SdSSdeMFFCeN0pQfJiIta3cuw6/o8RKYxWXb8jWeGJ/g1
zfPBl5Au5sfB9oJHLUISr3eQynOTXgQRf/9B65Q45isgsYRfn7euZI4XGLpVmRt/sj/mYMhT1fAu
kN87qkPJSmYZ95E82zLOTtSRb4I+eyebVv2HU65tXZ2L5JrplVf7iuIxRAzQwFwX+/1xGwwr86ug
A7YSYaLhXPSCffd2Plys9jxpMF8PaOe9VArWJwRHXj7C0t2lvLg6fpxQWLBDQvwypcoFYv2luKMP
9ijvG77EEhnXAzax9O2AmTIDq0lfYo1zMBZPQxymNlNDATtuwcxRGMFYExf5Ntp/yqXYUtOFIxKs
2pNly7ISNw2m/5x6FdJzqivzSONC7gIMqsjgnNKMh879ZiIG7fpu6/8xRmpWp7d6hiHzu/EQ/RJg
pK3Q5s6A/DP+yysIytf647ngp118dSpaJZH/Vyc+jDREFfEiA76nhXFdDcGecwDzChdpFkHjIXxf
wAN9R2SgcNDMP0KMg4MsqWoJdTZ0IwevxvACZVVentnKCzbKRFcbMnf+bnqS3qcSwDmeBlV2imTu
gvj6/D8of0aLU4uPw1FO8WE6kA8vha+hqdizOZBzDYgPIRJQL1d1TsKDugvEWMUk/VyyFG7BrcX1
GwBiUwDy8+5w/M/Zl2vI/5Bja46kkGWVjoIkSneY5aFb7FYZHXLLlKPns5CTMq3qHEWYxFRd0yM1
8rmKnBOXx2sb8pcUJvvu7wZtPi9HQ0nXNGJ9xuC4JPOmKz0S05k2NSt6lJ4ll1j/8gpoiQW7pxzP
yGP8LkqxNkILoF8ma5oWKx5Y41sFWmpjHvYEWNI3dgtYH1TZBKGVC0P9QvXjG1ImpcmyiRT/U8YG
K7GgD+GJVABjX7RGCuEFg/eZ1LeFUtLeTXUtxiUy3RkOWMmS7l6t6B0oMsj68sDxGTTCvHyoypOI
wGXj4VQI2H8yl89CQbAjSlj4C+pQVhGEegRaoRu6FRweAO64bMbx72KPU4rBNqB5BRDGbWE5Qdpp
ZxSJQwsEFeEodqnC0D7Ej1IUQrDoXloGqVp6aigNvCAzflDf0RfaH12cQ58XT7p1bDz8NBlb1CRV
ZpnQnlRH3J9OEdZSIyaGVyzxI7d5uB4pKET5HPONaDK/dwSuBDC5/26zdsvT0YX8/D/oQ7eig7iJ
IbJU06yBy+cLjzwt4f2VNLZRicBCFRIHe628mCrdNG6z539DTgr87lA1oRq/9zXBxpDfeUxQKZYO
h8pLP61ERFVW46fLmpcFKAvNoUuCt/QL/YV1Ge+tBMhQF4Hb4LgigzGY02I2hVTVo7VGCY2V03yI
1PQfNhpjFFY5JGSe1IMe9YJ8u+eImr45KN96a1/1gqbmciZSJah+ZTdXdepxuTuc0GNA0T0mfYvl
mx+fBRLyKs+1HwysxcTfwO7kNrzcj15kIriS0eQOfokbIj2JfecoIrNNS3vDfMaK10g6tPsMBVST
zYX6oA5pzUf7uVlzuWR9RJV1iukZjgK/sTvUf0x7Sm7N5XyRL1XP8oqLwcJTumaCUIuzUkCSnxXC
ETT12SZLZu1PRicHOvR9ArMJwZmizWPZA4Fondj5bolRgs+uwtWhub9AXdvdfw3uxKnnNXkiuFPP
2x2qpAGUlc+X2hhcXmj5drdNm8lXKHNSokILboL8UGZNpRfviX0ruNli6DM+gmAm8GAZhB5K9Prs
h/DDcELwjpfD3XuGVwP+ZpPVV2gfHKocMJhtbLizZaqa5D8lRWjtOurs+IgFl4lOIjkvxxoHSndz
z9MBjxwNFd1Mmv4sEdh9aKILXkIeBzVWj4sGpsgGKmJu3LB+rW7jommjj83JWMRNi6d78AfFY4jv
JoN1sOYDjhnT6GBQ+YPfDHkFa4h6ZF4pr4hHhsxppPpwl5hxuap699ZRlMp+1spJn9thOx6bfqx7
kdshD49ANvTo/owYAzpb02oQSDviwmSqY0W5AIR1CIiMf3moEtiHy669o/t/OZ0lbF+WlwBGF6Ki
eXfV9Y9uBHNcx0JXYfltbUQJ+gC+uvTvky3xaRVCyy4UDT8LiHkbEoDF6lJ4JF+UjyVKJFmiBDmT
8JD4KXAQjDMA8SVTM8k3YN4D8wqYc3raXsiQ2+NbFznIIkI5OISsGZ4MWmImMHOhKB7cL6YVLLAo
xdYFWzvcGy/gGxlivR3u8xEoyCV4Qhqv7t0YRbW9iv0LN+EjnPxV6K0c/I+za/3nKJXNFnExB/3c
BhlzlCPb+vewq4A8qL8nN1IwF/uIEKNYnkua3e2F7w2v3ZLtF+JqY2PaXkmgEONiGbeqBHNJdbyn
6yaclIR78Gxtb9bsyauxhQ7XUgORdz7Ogl+S3BbcXSlv++IDECjtzGGxsyqN39uVw/5MeG4RKWH1
k22E9y9fHB0IYvwTFySVbiduyq42m/JEjtR/4j2TMLnj6JqinN4DzugH1KNCz6iEbw8ZREZ30Vt/
pCWrMV1m8MMzMBuzWPTFzwSbQYLYEM6hSfIWefVbkEYfe4Hp4FeJwUnowHG0lPCjPwcLqs2rLjvI
wVx5fI9vRrkGKQGEOaFdbm4x8HMcoVSvPabyjtH7UbEhGSuzvS6ZaHXb4HFhvi8IVXpO6YRSmlB3
L47HR98XnHFwwSb6WVwkq1Xdj95Q/akQxk7vnWfmdhOlgn9MHIONHhl5W2cgnbzLvNwDjDw+Yc1w
DrHF70+Ot6QZK4m5BNIzsO7EXoLkHO3vvVGGNJSEani67B/xCZoNvJirSFlx9H7Mc+LxXzsm6Xp6
/s1meIVcE6sWy5AHuXhshWVZbkxxhWVPBszCH5P5I9Cgm7h/RCGH9Q86OChcHgPEiFFQaXsfR0wc
w9iehG9cXCrciJkNV+Gj34B/ugPth3wcCLOUdHkJGLSvsX48kTmpIPowQI7vGbqWhWIX7mjVmAhR
wMbOuQrk26P2A5FjW4vpN9ySxuwXr3afMmeN7DyxPmY8joXqde1kfTpLfm6XCnrC8ebWH2W23hhF
JPc396P+o7NvgWVMBjbDF7w4+aVPk2T3PpuIoXVDnJWmGApfysf5ug59Uj8kO82IlvNuKG9oVkO/
p/7VkOI8B9MF9FG5suZWrtgvS6une2iXCdEIOCw9XA7xqhEO83ydCSEXOFcuBQnkTycdU73gQCAg
ZRJ4cvBRsGknNHEL/r8MBRFcG0uWk6SEDe/xXyHESZZtP4SygiQIjbDUu3DG+1ehP9jGG5yS8Ytr
DK+vpD4x69b9T7r0U96dGKNiTBDcHiuuQYyJ4D+xH6Lx1MW0+Il9ixxFt0cr/yTbQ02nFxzV+Q9u
Q50KXFTCMuYF2hZGeu0q6AskaBOdh5ylVoTnCb7zlZxlmaYZ1s16A+STqgaC6sOoh1Em54xYjcCE
cJRnE15+5Fz/lbtW04C17BePXg5ijPVA8QMtuHdB70hLFQJb1mZ+exUZ3yJYO1z/sFnW3gmH7pZ/
Jz+zYAAuv2RWPZPEFtfZPGCZRotjymR4Ky+xqvt/ZF9iIpvAFPvaFLrBxnVz2zO9X24Q714RDmCw
hK/BOWNS0SxLgtqFqpbfaannQTUDEwZ/BdLJLb4YCeOArxaq66p+uZciqYAwzuVD4CuaassVO5of
KRWtvsyXQhfuFjws6On6RhOH2nv28eqy9S0kOE5nYFj4YU4cyDXmKI3sngA/JKzigGYQ2c/Nd3bK
Bd3fV07yQyx3RhICGDLt7QGWw2XdDVshCmlrmz7a+4CEk68nFAZoLNSp/8oMSkd5kMImRra5Btdu
ifOJImbDicvzQzJsYmpFQ8zf8HQFEko97UQm/fCXxkOwu+OiRlkkL54K9yXPE6iutQq1C609ntPk
IV4YMr1bl6pirsaCsTWh6twFDfVX+ta8eu05UWEUwgyLx/O2N/PuDRIvYzReC57nUvbeKaTAQD6w
SA4lOaB6Df0gnYfFOdA4O2HzEVFP7NiutuwbHUdrp1JdMOSdeRZhjkE/h+Qketm1t0XT0SYFUnsd
cZSG/TsYMgCYviE6Fn+SCcQGyjD4eKnkRQPGWBVlHPmV+3wxNovH2sN3X6msEtuskGg0dQGAd8YV
e2DwIQgoPX5riN36tTdbGB1tkzxG79i2C59eNMs8R+5hTeKsnTf9o4xcCS+o+OfzzSsFNDtknsbn
HS+RRJaOEKIaVCHsycEQEzQdlbV/c0mnF8dzkimNZ5lw2Te77TtfQK6b+SZzK8POczNgFGteYlca
iIjB43drgPxiP4jEBVPZwlyNSAVVZvD/103F64TYZ0i93xhesZXGg11sAmPiGfHDeOZ/n45fMZwm
NHwqleZV/PAZM/2VgZgsHZ8BtEMCBUZzp1fLewPNHFCEyYTE13cX3Xwa5+Vfpn/ypGdU9diLtC0B
+w7Z9aiEg9wjeRup071SviGO5mqvulboXu71EuXg6O4mAl0BwiPv4vSXUJVarxS74WYAF2uFm2tD
6hxXe73WQHthyIjfnq4eggx/zjpvcJd1cUBwRxqWzmFRGJh8L/Y1Spdz8u1j0Knj0i5swww53yQj
6qdf/+MgFWiLxJFo10Aj1Q2CDwXdUcdzQrsnBwnvIkw+VzF4vGuMDrIxxydGhl1KGuw/cieeNYVo
FAMCEjzkMwdXIdZsfFE0Pc22JnzSUCfhXcvc1yW6zgANYClIHafNfnenjrV55IQ4QDI2tNXD2LYX
UvaBH47j+02MNSilcQ0H/nGH3qRk9qNHanvFv2T9v2gEeITcK9MD+QSJfMOwBp+MBBuvtBlJuENr
/n5+iK6BRvRKxqWPiLQMRlPcfu5iKVb1urtY8eQ3nG15QwBn3ahKbCo19roCItibdzbYwoRxdGQt
ygvJmBuZJ+X1Hu0aucm34jiJPgtwdJmWa4hrlXJuHXEZOkwbyiHespT4N9vn0LjnmoIPBhKbfi3W
3IkaJ1fsDf/wU3r/NTNSXS8v0M2xBCRh2XJq3BvGXRpgxMWSAbeJKdji8zsCoOQszzfguLQcAFcq
nuKosQUZgPxxudrvtoVF/Cskfmod/yHdITkzyANCYz1quruEgNaFgz3YHzHCYoxBRRsrqd6T7JC3
ZHXvnr2QUfor+ytvjqyUYICYtDapticqC6wZz65ZHSHjf5adK8K/B5QJMI330VFNcYbrhCRZ6fmw
UH0ICvJg4sBif33vOB0RkxdtrEdPURkFJz5u8LWUJwEV9sdh4dAVeXQzuVMEX3fkiN0aeoDufC/Q
nGUkJtl8F/V9/PZRm5e+yIfTDeua7KUPxTtPHoQADaiRWRt9I3pXn0DBR6G+edrooeQ1qi0DHGYi
uxbhZ2DOspC+WHGH9xap1APCEDqn2bghbh+/m66TSm+bQMaWvOh+axufeq0FPGbbpl8KxVonqsQR
0HkdS1UNqsAttmnV3jktzYsg6f+WsJW4Z6iMq6Ri5/q7VtRjiCApTFA9Pur+Rih/OGpcQ1a9FpG1
tD/IhRPVgzrhS55B3QQg6w+rwB/vkM8jr1vaufR7PtYZ1c9VafgcdJ/xAZNMVQhgoY69xrhpm+10
rZ/sInui0OqdozKtJyXIp5Nbu1DMefhIncib0b7ZFRD+6b18Q5Lr346tXZk8L2OA6CiQqJYxf9AM
An31y1x4XdQ0ntW5en110nKqVi7ds+Qq+EyyWo+8whakfgsJ3ELVJqXx9ClmzrW+ZH0qa7XrhuAq
gOSPGHCxqpEl9U+LSi9pCpwL0VmQobwunNi0869ZEwv1PMaAdauxpPbTQVcrKIpubCQYAzaG2MHb
6EnwbK0+Yk/iNB3KOQSQrNsOSC1x2O32wJqkp6818/Hv2dvre8916EH3S8f59tbzh668/pL9Ti61
nKRYhtjA67LHyXdOIhqXAZNEiqQ+E34AR4l2h3o+N1dZPJi6pHOWSXbBv17po3ja8Hdl+kr07Prs
MQePPMZMSnLtnygABlMkklGzGrm1nn803SC+9gryMFm7LdvXFMZJATXLzIf4KvizmpZvZTsN7/zE
27Xenm8yDflb4hew2Dem9AwnKQEDgrTHfxnFyPNUE6U9bldaCjrOQx54K9aZHxv9J/d9w46pzdew
gj7Y4bcEUyWFrCQOmk2IaPyLNpUToftjy8/rPWttIv6/PBvWF/wJq9TpyhDq4vL57yuAMqqDdVrR
7s/30ujk2H1jbTgjdN4o70PjXXkKbJ9z8KM+euTL5Yo9tEWK51fNQmnoOdPq17QiKPHJKfzI3DU2
V0z4Jk/EpqUl7OGV706Mfe0Ps+nlsZsdTf9UKT4yQcdt471dyxhGD9JJ48aspxD07PZYZZBv2Qky
2RBmmIkKNrAqAbUr+F+vZ9yNoEZZHHZWmQtI8x0SjBIBzoPZ/r5nkBKHkx0xMALjFerBln/pdWOj
lrMGLf7yh+d6/Dl2HWsJLHHWDS4O+Kwfy3HV2AHPYhU3wglqo1/pFN4pxouWmlmTVn3DwlMBioi9
zSOOLGMlM2ZDp8d2YCXuKuWDyp5hPf0SK5C2bFwfCu2myL5oWFWy/RXeRKv+Ar7HjzZ1gk84ZtwM
nCGudrpoKQVw6HiToAOy71cMnd5xUtAIJuXN91+UarpB4IHftYO4uRHNk5gilBhTVNnGP25mneDf
NjAlEcFRevHeAn27pPb50sjxsZpBJz9qMeo6TA1o2VBIsjN5Jl5gnB5rQbElDbW6yn4X5lHyUNwN
z5rHonwnvTY4wDYda6q/XhRiX8P7J3P4jZGdWTsciaiUvCM7mNeLLgnT49JoobsqtFKONN9C8JVh
q9lU00lJjHqgB9Rh2bTNZuRz2KTwrW+cT44YfdMRcj4aHh6EJUFBHEmbjqBKvQrhyIEZck5v/mSA
J/ocY6txk4/DFUOiqFFqi3iiTSCeE77rHhStAuWEskqCC8YU5N1C2lSANQKWeYIemVEdhJMy5I5M
Iyl5zp/baTlBc+igxl8BA1flOqD9M1lN6uGhtcCLAe6cpm4gt0ICQZTHq7vTdJqK3T/D+u3wTO0j
yZYEhbOh1LBdr7+5uFSbVQj3Z2zkJLDb1hqEBQ8QdDN+iNHt3UwjKVQ3OiUkBml0G9DDi3XRL357
71y0tdnfCcHyilk4tlHaa7Q2eCvPC5mZdqwCvbhD8bTm3g3JKcM9RP2r+bhBRfTAzl0GkhHB+H4z
w2KO4ldPruqqBeL91a3Z3A+kaoBTdnQV0T263wnEurhG4aN9E0khlRoF8G1848DZ6GvdZQN5sE/S
tJ40pu26kO2fPc7bcoXZ2umiR3FQ1Pmgcq402riAGwvbsnJD1tfVguovLS5B6+k/qoIrpjH4Kwvl
clhsv8YKRyRP3dXdmpmfs0Hjdy0dNW+3KrBVDL1+8xglkhzH1GIrRixcLAXpNdMwUzzo6BzEgzVm
KlFQvJp3TFY3xr6wh4+w1hrdLap62PhcRPmiiLEjh+lzwJnwG67QuJS4ZXn3GYu42iOPi4OZ1OPF
G7LgVcJVahxglz9x2dXLeHrW6qoMlGnjN5hy1DnWOY3LbUyzT0tYJenbrfU2TIrrqod0TMENH7H7
3vaRayh0uU08NyICB5V54+xxynJ2pK0UHSEJXy2efSY+7pEukcW7auwd76UJda+Z8ktRb05Sxas6
Q0nM4mTZIG5SsMDQpfAytCqsI194ozdXqKq2df5Mok4tvM436yQ9afyQwstVzl8Qzhk939wq5C7A
rVRdYu4kukxZmwYVwFkpK3A87G2iJxEA1WF3ryFBf84H2Ca++Qlw3mooDmLdwGAMMNViJHLYRkGY
avQdqRTv/AZhHS5n13cg/aABXgvDjExw5Ock0i7y+dQ2ZBMv0TA4/QLM02YEfzBvf6iwyoLfYWHA
t/gX6AEoXzuw1dw/26fC4HnrQr31TN5h38gkrCcl0XIC9bA/GxSdobNlrf2MQF5AC/6Lc2Jgptfe
c/riAOmnKT05gzUGiITwutrrHzcfr1eBf2LDRIg5fxc+GBnWFyexWdgWo5+UQ8d1i/KbDCxtLZk6
/vMBx9Y2DHQn57SDep+CmwJzAhIgsPz0WaCrM+Q5LwKcZ0MUhL3wj+qN/yJGAPXN0423svR7JHp5
ys7MzjFFd3gwm+eSAeCgyVXHuc/HOc5sRUWGYDdH4YtO51Djst7xSBGipkEBlX441ImWQBWjFygD
nkH5/ULyI+7mDVv/sbsYNgY1MZhCQTmrCwT2KtNyC/oDVupXOErZdaZlU13gdNcwRBA+Sq4ToOm1
/J+dWsEy6PoPCsGE++wxQezgFKRDxuAdAK5o7Skk/l3Z3HhJQ6IWZSW0Q8qm1/I1R3QjDbDGMTuA
3jT6BOoW7AeRTGGEQ9zXiU+4f2d64e7wS/3eaH14xy4VWapyFSStqrALoPdIz1YzqKpMJuXTsQu5
ZxokXPW79QEISKWMrt6+Jqqyhm5HZEy6CnfMx61VYv/EbpdpuLWOsjPSPEQto/G9Pj7s7M9gXIL9
aYkEBJESyuzDhWBmV8FbvxNbEF3rXlXEW6fCbu53CqqdV7HtWTUp+3qiBB9R0I7JqcnAwStIdEXr
rJgoGGOBpGzPOy0yEvvLewH0fFLrjx+FcoZxCaFlIDgr7Rr3IdSlJV7ELnWK9kdk9nZYLhv0zqlx
N3AC6iThKV3nh9KOymb7glkPBINjc0gUskfWDyNmXXfxanJcdLKWR/s+cCCijwJE7kHRNhrhnKEa
E7BO41I9Yk+kJVleneTPYJd1qGao99VksgfPdtwURy44sk6HYm5jpRRD9aNI3Xr/3s2ALgvzP1y0
YIEuxoH0GwfzPU0MbUERyKAcmYAAcSaVOPWJUmADa1WxJQw/61DQz0/3p1KsoTjBNXVEkh/Gaagd
OfuMghVQcWZJZCiEM8nmg3igd+C8M3GD2zgOxBo4xD9IuooyruIxCNZnD2tJY/0HwY9a3pdLdAkF
AohD55EUdhTJF1X+TO1azfNA/ZZRU7j+Lj0Nvy+U+nMyOtc1zXZCQLPSiQqRstDh8Dy9Yaq3ehXL
54zripup8h4mqAXuHJczjwlNt8cW19wn4kE4M9RzVADcH5rGkYZezu0eWYp7dk6e3LWSfv121Fn8
hZXWAVCfai5D3X50a3iZ03US721FGxVbw8uyC6PUvpIoRF1mKcCB0zaC0ekOFBS91//h38E54p5A
FC7YhE1mv+P0vKRjMzPSN4q6VdUrUgLInzoIGj4h4ufMC2ClbJgwdXhTzgDJYA1vjfAxsXyKPYbo
VGwPJmxIyNwbxhZh8DyZ4r5O7sNkRLldD9a8xatlyw9Z8AHGmiRuFFD2Ua4DomhghmPSqDUZX5jG
YfpsZTiursvol0RjZ4LjEXl2J+AWfFKDAUv0TNhS75+6kZcfBJ3XWF4ywp/39sYKk0cTrw0kSe4T
ylmxDfSHnOwWCkFgQpRNuxJNqPdce2mWApPCQ0X7544cL1kzs1uAb2+MA70ViuhgU0sHPvC6F0qm
OqMz98iPLH5ydRuZYmWPA6my1yKO86/M3HoqEos0UkH4hTs6McvSmtRWuwBfGr6hqhwTfEosQjNL
riRXi7XiytFj70X4lGX78SYeQL1Z4XaJT1X5SJZ0CxA64Zq7Fh1wDq5PI3Hp1Rmtr77OhHAA3doA
V+EbfoSi7IeKd3gxuw1kg9y/p/rp7PeHOkgV+cWTqZiiHb098VWHMp7Typ2qFvH2mrVlzyR2tByA
shEcMD/5nL1OH1rYPibNfRVoVBjnQhuNQuugGk7QjM41pMMNN+hL2MpkUHeW2fPUkLIh9dwedirK
r2IwrhbR2ccWxq33WUYya+MYcRif5KDxFu6dgfaGZya4W77fLnh3y2fRWAq+S83V7j6gr1ao3nYI
2OLf/lMjIQ/RSnc6zoO3XJ0DfzZCwSNZ+jQMPFOK5w86e6lOKDRjUGutCtGwSscbT8XhA/zq/xW8
+fj1+6TaJA85oyiIHrIUrcuDQdAI2Al5KQxYbFmkj/fBetS2xQzGtVOWjbbpNAO7WHOVAdknUgmc
w/dJPaMcZvGufpGbPpRZtVXh5ZNcxFwoHNLRE4PA4R8wgbb15ul7tnJu4rNQsnDyQkLwU8ic/FD1
clbbUpT75GJnO0utl6jKlbwAzfPShbh7RhURkDeX4hwAke/OlJ1uwaej04MlfSHDTFs4VlOzdnY1
A2ebG5a9Mx5e/YZ12zdf6kkl+XdyEfsTesCGQveJ/VVhM5Kw9DpGanz5z/HWBkMwYH2A2OPT9EmX
r0zQt3wWWi9Sb+nFcj71Nv9/Gii10UCJXL4Nyi9g75IXZREM0x6gAV1krIYsDt6ltpzc2k3V3NkB
NYoZ2IkAInSrM9ES6srcJh1HLqXUhee79KhRSdyaNgtXx0bO/M6W+236AN+300zZf++cKjPmzXE7
7JkN39G33TvxUNRl60ya/ueMsHoUJamSCiJImZBoduK9qIkt4+WDP1r5cXck+qd1wrqPm1UUoOwd
0a7eDP7j0ucDfkR1KrXHs7KKkohWQ88WkPG4jWArAaanG/8J5P6uwXZWgjf3kLE1VTWdEnCLNJQR
3lUE9wXRYaoONmBjgenQIGY6GsJhdkT/jxTaiBal1Cd5uhxrd+IYZd4NtHiLHh2XEaG/gyy+N5zs
ZMBlITilzv5TQR/pOrclJ7asz3xoOKUOwvn41WwDazH+XrfAbbwvCu0c+VDbK9iqNi794tpNU169
Jxh3oHvYf+ca5ygbTVY/og97JGrwPLfsUQXyNUJ2jOnQj+X1v4Cz0/NyaBQAugqQy3peQMdoql7a
uTB2EY7BZ4npfW/092LssRSuDjdlyPF6ddPWUBQtGKRwW3FX55gR3C6odWRMZG4717aZw0xU4Q48
qH5vQTfrdjXSbBn7JzJB1E1Z/xQfLmnUHKd5/fqoarAz4Zo+1e/KfiVIuwlDCwk6FTIBh6cqyHtp
FSSd9EuIKQEYXGicu+1aVQuvBZPxoZwpgWnK4SQDWz6a0ZXMUkFsPHrG/u8ttLDKfsm8mGnAGbVC
tYS4noADt3uCPC51B0/o7o5BQbvEc7VbwCvUm6Aw3HhvFPXg17gzPFBZXgVQ32EBo/nciTOPTIxy
xSElnrsbhcY95ZM9nYsQ+V3KhUra7pso4JoCjeGl6bNHGcWWX3xpDOFjJBGm/OCpi164PTGvnVs2
KHillhYUavWGIjjftQrzHY+e4Op3FGaw7taop8hmbTfCX6gdo2+QCGDI0vzIGhlolDyYRoSheMi3
BjBl8MJFSuM5xwleylTVKlIGKublZkc+odVNbGa+79b8jLGv87UkeD8L4z8u31L4CXG/+WGxnLZL
HKL3P2v4wndGNf2XDRMarHZpw+NckQgaqNAeuMUHxY0ju/dvDupdSwlM/nd3DgpHkUnV6a4S3SkK
99R8mTtiK5BLjhccTgdchUi/5xBuqsd83kHGok5Q+qGYyLCCRvHCKCarPnpwBnKkscMnD/1Wj5M9
EZYq4cXdl70b3QVxkB3XlNNpduR8KzL4yrhAH4xaF6OBupACQBX8wMrK6aKWiiHQL6n2qDSWwJP4
HhGtR6TO1By81IgVqE22v7+hnBhIoe8/0GW3oI8SInSVhNLM/TZ7sk3qynESzBMLHes85wHxNxPa
Ln3LqK0UffSN8M5Xbx4xpM7Ix4NgMLRqqcBgyB1NfNWRlWjPB4FjFIguatLLx4KmeGJ90gF28A5c
rNUWlHfQnyNsyJOVaZdTGNWh0UmJuDnvzauoItdLNSPxdc33QekjM+4J3kYnRcWjVObok+cSR69+
69UDIYxrlJr0wbd1gxycy2NNYwOZ5z13QbdS3l7CHZjKBjHL2gdwaFRGJErfgw4LZZBX7U0dPRmg
R/s4fTbfo4SZvtfln5jcH67HGCEh4Cc/GnyYTwbIpI1y3C1m62e4wbX1Snh5jHtH07rB1KRzembw
gBw9/9rvg6NMK9iJcNrjMUnLU1r9UCkB6mh5WYoATL5CECIAOhYhLQPDid9FGT6R56vmZJkdOKhN
kcihnC3Uzaw0YWIj81hH5b/vaDojHTN6/8e4jW7dFeBDbYdny3CeAmtVpeMylWFUbojubGTVTNey
cs5esgn4tHZee6oYNAW5wGYSTF6foXhbdg3qNoBuqQ/bNFwrZrJ/cFk0Pe9JDH5zJNEBY4Tp46S6
F8OdHUqiV2GH2kssf0pbMVTPPghnCkfwzf8OlkItCZE5UiD9u6EZ7FljmC2JA3qZldH3BdH0OX6w
zrM5Hn6ln2SIP2OeEGXdBQRDK28/xTyao/xQWXk8jj0Zp0mBdBXcjCYk82rka2pqJBjxe8eoy8if
VQs5eRdNh8IxIi1RaHa0E7lPyKpRtbwaQyZaqkaOLfo3XxBjMRE9feQ6DqVAZMhnqNqLisbNaq03
1QBKB1SNOUCWpee2eXjPa2sBA8+tqHQIfg2X71c6dxe7vkP67ErmHqHyfwC9wpq/2as/g2jZnrHo
FHQRH8EB8iw/gmrqmlWGrwmsWKt/XzOW+Z0neGCU/DHWX7AaGFdN7997SDlzyWAgqSrQoN2qBeYe
owCLfX0VdnCvEfdt0MNF227gODBY/Do9PkCJKm0Ula7PqHDcQAOzPlRpdSLducQlrmCKSLiD9KgN
Fwn+ElD7llX0B1tvO5FH+w1bT8EbMhcGjtXKbI1xGTt5lKnHwW/r/d+dSUziO75EWwA7TxUhhEq0
wMoJctHtAgqaiqRKtUyegqVF64go2mFnqnnnY61ky8wOnUEMeIEuf6ad2vYj8kuisQbGu3ktHqg3
z3C2O7QIfIvQmicVSwr7EJBgZiy6xTAGPLKsRGaGEGlS3iIosA281jYslyeLZq2YuAVS8ly2rFd+
CxhbNDVTuLMVAqcGu6AXjNag/G21Oq9VxgZiEdorpSH5LROkXO1McVTtZNcyZ2UipULDxvw8CzKv
+wjjq6wSw3qFt9tMxYVE0/cbS84l+WS/9Fo4sFGEgucEO8nfiusB5tw3VSJBVZLkOc31j3WJO+d9
nr2ZtAAmVHbbqOGRM0OQ/GBQFwwVumwO5N7UChpXCJPFCoE6MPs5C+10ASTePF3re0DRv4Dhj/an
EBVF6QKVOhcuqLGQoE2Jx/nXMQha+X7PItkwx30p5z6x5U9Lr6KbcSXt3qPluiZcXqcdv//uqt0K
YtgB3LLD5e0k8ogv/8m6AnEZ/x7pYGMuPcr1o8YtO5ue/R3d04M4P0X8i5lF1CAZ6XO2zuHO0h3m
6Bzegqfz8d/0tOei9jMtYOeIDVPE27rfeKUioaL2vHwrCHtnQrQavomOBJ5CNDJeD0pSgYX3jvuI
Toxbr0m3ZwTW8W4DAr2SNGUXjMKRSu2bFipvGyF9aJ2O+qoZr0IaVFbRfx7FGsH5jPXpkqxFPL+k
FzL9uQGhZCsv+dCe6crx66OrBgWC58+7lCHZo8BcJtNsRf1pspQAB7Pm6He7x5ANSREd/SThxNnc
8RRVe41tQwWg2HRRgFkkkIx8Hiz851Qwix/qmg6FyUzSrcvMAj31kxq/NP3RsGnLJlog1XCpOh/k
6HMyk+EjBsh+/xDJFv/gPEdpO4QNhtntAvs1yPw4aGt9W2GLu0z4rk0zLIlZ9ODziyVmipkDv4eW
Yfy0pcJxF3coy2KlJRKrsYaEXbQ/rHdXSp0+qUUkSjhuj/+26ZM5C1ejP7IZkzA7ZILMVoFGTpoW
pFwjLDDzAfEqyrIyxs1iYUcgLajPdNz54YXr/Je+kaoL/jCOXyxWu01owCajhUnzyi/jBBS3zqIH
t/EtwcNv6bVKi2+vfj4yQDNKYHd1QWfwm7Pz78Zy3XqENTyypDYjvs9km2tUZUXl7zrvm9stz0Bm
mn9R6eoYll9QF99kDC+BbMXFSi5oaPmsPI+19hQc1P2tlSe3fPToYgoEDK5hkQVjOvPTErDbHjGy
3dAaeujWcqSwW7X9TamiVA1CbddLlMKjSIAggBMTiLLr1xFztuz+ZaHAW77OJL7WwqNpT0nCueDE
ou63hVi0o3t2pWcJjmEv3TfYeszlRUkzCPAMSjVt16mwtKX5fWer17QCrQ1L5ix8ycxEIEa+dCQH
SGyfr1t0vjquzI/HE36IUhidsdHTaL51LAW9WqD5AlmFC8J+9Nhm6YPbWgEwzQfHby4D48Urx/8f
QCy2DDpPYdgKLWv9KE/CdK5ggiGZGtCA0Qg16FbEmYBA9gIu8HIu1y8FcjuAujThw+9BB82KJt1l
tGoXLRNH2kTkhuFB03v9I2YPmzjktaYbcNy4ym87DUyLRA6vqkP+YFbsh+thS0ETMZp1ffqjznn3
4gT1y5YYzb6GtukYH0i3G6/n6bSw2m8YtoT9ell3RBkvncY42AKYs39k5xQocaOjxO1B7JgnJuGP
oFufDitw3WzmcBxUVIHh5B6Os7YJ6/pMatAXhyZrsqGcdpvhIdI1UcxAMuCyTmmQfkxPCPKhzRCs
u/rsLw8GAnUexWWORVxEipApe/6O1KAxRbfN9xWdrDb8Nb/5w9Vfmot3i+Ku4/CjoV/9ahRUuS1J
s/T7XDzlOROSuwwGjoY/HmsNLZOKoYb0uOlpu1pJ42GEslBcM3JEFhmsTRsLmvoKLGExH5SBwADG
dldfiL6U8yRbuTPNqeDGH5AyzmLD64FVI/dLfPnyrD6UqE0CL6nPnbVW1PbJE01AMRONok7WF+jx
FerR1AYlK/1M9ApSR5uysU+3GsK24hwrJYwfcicPFSVsSJZf4PkrOldEqKIsW3RDqp2Q2/mm3P52
zskjVPBW+lFbYkwu6Z4N9OB5SQrb7keHvfaRcoAPsfP+FfodU00mAfDt4R5SKvLuLDUmve/q5X0v
7AMB1PjRsMOVs9F6kccfAzZg3YDPEww6D3o6YIW8en4zrGDTH6FYpXou/UaysLdmgGGBG07OTSsE
tMBhkzsnX6LKqcCq3EH1/pJ11NSEGh0qt4esuwTU5Zz0A0IDvJ5Yl7e817TmNImJAM7qH6lYtGvm
tFWKGYTigj/WlC0P197VbHNzJJpEw4wXxY8zQuepAfKRPhzGGUw+eoZNMP1bZMh0g7xCecOKf1dY
W+Ot/t8NZxPWFA5Pi2WvE2c7g9o+y1rIhUJz03cabJO2441wGhI98QQtm3oxKl+M+t6d96dM60fa
FHFKJzIjex6sJfJlimlJEyhrbOJAdF36TjNj6Xt4NZ2lqDDysv7RH/S9NP6qsGEt0MEPnNDNMR7T
krSn6RgjfOplwOjchmy2eeJfyeJve+oOHYzu6SvFWzSkAWovJgnkqICuyf83DodAPBeXBCoOyTXa
nyZrv0iyS5sGb3wL9b6HfmqOoIxSRMoZiDgzPn36OKaqWrFaFkB0dfWMO86ZfAWK0eHa8+hvYL63
MvBhlFd8kFB59/hF2MOiSumbYTwtxxoZ+pTtHLgtWp44iqbCS8q+hjP067Pl3X5aP4L348p0rzWn
2sJWiIhfKQQzC5KPbt6+ivyIIA6+oIi7jhf3Pu54KQcxfMmNDChP3Zq0rqM+pqrI/B7o+at4c49p
u7lKIUWoFmFeXM6udKlpAhZGIrPXjzlqHjmRhBE9rHY9LJiPsw8Lyg56K9bu0ny4rIutbrOsY6XE
KG8mCSMnZPD6tGZwRvi0lSSsClaZ+pIcwxD1OMDczwDoWYN59etYK4alz144C9TV4V4rom98njrM
O6hSIMVl22aodxNPJ2SFafrBtgQJThhzUkXCrpv9Pvr57Jzvn9ehVBd0gAENjyuRIQM/Cc0AJoRa
eK4Wjv6kaA0dLRRrbFOD7+a7M4u8Ic8F/c4R+m1GuASjdQFsCOE8CXGEtBIwcI171cD+ZStYbz9s
ZZZvOk6Y0gFjjSXRpWCRRurBmfDcIVfT8rgSt/LMshRMiFMiviQ99ckohaYZyebQOcCvUUPVGN7o
2xVOpN9fnHwHyrvfXWUqaiesqyNSNiTHekXlsAFcKMtcl3s/yvp445/55tFrMQ8IR9cMTxyDAI4a
qEajlP2ext9SXl63UUYwGGBI1DtlJpYyGQJ5kfT/8aB6IO3nkAsMJ1+ZNwDoBs/k2/DGWPZx8AFJ
7qCZSo2JjoXEnQSnqVvP7KzC1ZDR7/tJT1eABOdUdrYTyCWfxrYS32F/pJ6q572JRGZd9TNbGdDJ
YfMOaOBjZUR05lZISOjRLwqCxdQPgZhtFfDMVaqn38fkYWspQjXl6StU6G7gBvhk35CCXDRdAzBv
Yckva3fPf7U2lKDyFJdoGQ64l5QAGHeMP4jAsBp8Ug8afqtPhQuU5YuXCgVAkRMc9UnMf6h48CH4
Dshz0hg/Pq6rTMwfdBL1MtB5DRe41J8rF5h1bumSGlc+gbzGoQRNorxpLlhYw3tkxuKAJr2ETc27
Pjirg+h1UrWWmExYYDRcW/NeYktCuxJSxWUofS3bAxQQKsp9qC9YEyl+G0PZpOKp12K09kQK+eK6
YPM/sXatOfttLg8f0FnqM5teecELKVa4rxbd4LP49T6SZlAbozr8NW/nZLe3IfRtYpdKk4fSOPt5
keD/irQyfuQePhzWe5ThoepXfo5O1E02BHCaA1aqdDvKbvB0uvYMtMpLxeMAO0+RuVSynexf559C
aZcM2DOb4GLFTqtRLe8ZpP+w4eGMLZi6zZvyxR3dpmKujBZ4vu5Uhtib4Q4JZfO+C5F8URKwQdPQ
pRGEkwcUWLjOYUbWdi4VVs2MEFyXelO6Nw4u10WU9isxznzVRZ8SxK+83Y7ESR77VuI7HHv/LfvF
F547K5+hDMeNY6RNytx2BqRNUAL2jS9XblzLDnAeik0/9jsp7QSlVVltiS+0ShrvkfBR4R9L7qId
K09IJULBSLOR5ZSl6wvg9GKmxWVn2XroYn/Z7J1O+BTY7kJDLfA9Wm/bjNXEE0G6di7Nls9jPnQF
kCHFipWSf5GYLNq4VgTcHA3Pw2olu4EI4U0LXBE07AsLVm3BoaQ+54G2mRO+ZOiy7N7RwYJCdQdO
SnK6MLdCjxPXID1wtzByhh9ZarordPVmMQ6Hy/b/lvHpUMRBI2c0J6DXajfM0IFVpnoBqP2wQ33o
39tQiD5cFaPGu9Htkeb1Gl04A2h2ixUMKo0Jvmte7JI5kYwX9urykJDnCbaLsE6kA/lmQPHh2h3L
Y5QTP8vwVzNHfAh8LHqyjpOdJ1jM2PU7Bgpy8yi21IwrH0RCV1B58YFKUexTgKqBwhnWieFpJt8A
vPMUvKWOeMtxAImChwAUHiDO+wtzPMCe421jnuT4cAwZ05Lxpl6CqZGYFlm3GShQIfot0ykoJBgg
BeQs2r3S5qV0KzWGs1THDoz2NcelZy4Mgvypg8/Z0JmiX5iEoDdWAEZbBSS3Ul+FmSb9KqNA7X0V
tlOU9d8Tju8J3fs/PE267GKVdZywpe5d57DeXF/FGWHaz0oXUzeut8+lwfdXS0vJCOYdiWyzvysd
//bPaktOqDJRl19AfWNaAqLO/hSAnWjtIJVy+f9ahsaU2J0BHGnavUECDpAO0OwpRnJ6PzGJXTgQ
qR8/FZQSf94nSdSsK66OPGsAEcfPkps4Qr/kKHrFwdRx53npxx/BqUdF9J6Sks7ceVTkYNvLmObK
MgvgKO836/q2fzM5cnYwpjmR+eayq6YU3LWUmlsbttmjHft2v7RbDuOyRSLY+a4fJ6MZvTMTxgI/
+SeLEk415MoTVuzlfSPNhnz4ral3jXmHoWLg9vlSFgV5bk4hKE5lA8OcNxJGTJ5IgbjLB7UDC9qV
VXb5GqG/K4ybcxra+hvD2JcJoFPGSeJcimmxgx4XnGeBu78sQnzMaUxJB/hnTuy4D3PT4HIrcJwv
gE4/VnOZqo2uVJOC4yWtDMQcb/u/kkIjGcoI6qDW0H1B7mQUMRG1/TwI7eHWc3XQSS9pJb+VJ/cn
2FkwEdNSB/9S//GHqN0GD2W7NTa9D3q9E+t+3b83IW1HuWglPi9iy3AyBPe1YwqgqQk0ky7kNY7K
j8+dvtWeWFWf7dsEJ+22uDyVndyrOC+OM60cfnngJMH9Z4pFtiBSxGNBHy8AAojj1qKXfoDXXANr
u+Qte9Ko1rzeNs3GkrkVunkO47Iw1Ed2aLlGvmCE/tWYM1iCelZUCojHa2QQtmQRJ/2itDHzR00s
XaM+5RfcTQGnV6Prxr8g1FcZzoiR3Bz1H2mBRhYXoQT5GnW8hZ5t4fpiI3uS0wK0toaq7qRHVg3O
alUq5WWVc089yBpK8MBTWPG5eStkEqeK8lNN1PqZfvsUj8TmdxLTFa38cX7CAVdqg05Gs+bk8/Qd
tPHjGJiKqB+GeSHPb6p5FJ6DqzX4zhiswanoa6uLmNadkevi9vmcI5H5JbZngEjhWEoVHtibD7+O
PFCnrw2VJpiaz7PugTSgNVRJut15G8Crua2tLpEjxZF1eFJ10XYztkGPTkaYeEMOSP6XPFLdKS8c
BmUOgVDoEXIQkkOhctRgEb1lyJi7LjQSt0PbioHuOQtLJpYnsyDCpC8Z9Hw1NEQq1VZv1VPZDmOQ
UNZNKEbmNvKS5GJXdDIdaTozxavBcZvL0sp+IYxQ2NaS+BfyRCMniZIkybPUlW8y/OzFANYAzKNR
yVl9tUD+KhY+s7IPqBcnZfJBjEth7x8TezGiwwbTlBO+AJ8YB7ew21htlDdcfQz7jJ8fGmawD/3k
qLH34ahXSRQnml1bV3umwcDclFMiD8F3QIJ9qUdMvlkcxzuyXvtm6KEg5Eqvzbdp40UG+Rw1cHu0
Crh8cwkB1oi/Zm1Yw7Z8yYS20aeG7DgkOSmt+87ggfCiFa+VVUvGCFc3OIROCWWAS6NOW85J1h8l
9OMOGPD0SanBr3UytIwIBpORdV9Tzufl+M80GKguOichLe41Wg09HoW7Oxyea5TLTSy/s3xTKZTF
tRnuUO4dOsOKHXD+QfP7fZ6kYKZTb3SlNIuSlKHix0ybLWhjUTm1JjJYvpY17A4Qe6xlib+oZjIN
fdM0WCM4wbODVKl8Zz06GwWJtBBh4+Uvm9FlD/lkxmkuygTZp5Lm+4IvITpUaeZRrYkNSKqPmMNU
nUP+uSlYYuHtQB5T6RPZp8FQwwKUFuJWi2PeKHlbq2xq58A5slotMAk1Wb/VTnZKg9Enr7kbEiz0
rM1pBQ/cPAkDMq+wGSIobVcddsAQaN3n4f41ssrr0Y1rDpH/RdnG5Q4326fcgM3BlaVV6ywzi8zK
955UPr0/ke/P6VXEM3qIhcMCNoBO5ctpMvprn9Vn7K/1Og/T3EhGwdU+WuAuFaLmhJRXyHfyRB0o
um/Uh4VsZHKyDJzAed7qR9XmVHO0+y4EXYK0TGG1uK+ggC9BBywOfBBXIlA8zPfSI2IgNcC2gqp7
C5VjzJYMfSou+yGgGBRdcc2vNEykc1f0/99UT6vGH3nlcAY8/WgHiPAX3biFANNKju2RrUxvdTzo
2bCrw70H2Nbs7DlM8Qzfis2bm8DXGcB58nRUBHEv/LsM2tU9Uh0QIJEfJ2+RunSXORAKMKXpOIBG
6E+hbnbcdGetUOoLAWB3s206MRJVddxfNRQHEUDIuXJWt7A83JFUlu2/AEQq/DmgksY2+cXmJpnr
mDru2p21Ob+kllciom3d1ZvQufMjTUtKQ7Q5l7LtAXoPla2ZNfvfgTeJmbW2O0L4KrjN0HT0q4AD
a8vJTpt/8SpjIP2YwBZZut64qmxOw3L/2xuHGxondIQKIfmA3dzKbVeoxKdQJS+N+q//imPK4dtT
C4wnFvYc2Yca8oMCfwtgfQ8rB++m5QDEVgpQX6qMFQRkscHtLePKj60Wle/fjxdI5tAQF7yZHWH6
lGrub8ntbioVTlFMkrXwpLLZgLzspdsva7xy9ZlIpQFaStoi/FVbOJuRofFkY3g7tdY4rZZUtUWO
nZmRdlTVXMVJ37O7oPjjUCZi13ShT/P4lOsSY9XY2AxKsou1J5WJckyTLp4Ih5xTOpsNu64xKi90
GSTMPhNyKQM07ZIVYEwMOd1otzgWDT2+t3Rh4XICPn1xg/WYexArhVPepQR/DW8aGjbBdqFyRymv
HfIAmJYqGoAgLN5QJFF9coRUGvIM1P7u3/RYAnEA8/SPgI1J2Tx44kI6uC+rGxqkrtDJh/S3sOz3
rdjmu5QZohdzH6FIFE7Id9cBT71OJqFeAz8n/d2p4AFk/N8FppIta4lWdQG6ZvkPQxYHslbpiNeP
xKUJrlF3/DBkyndDgjMX3SC9ZvnV4DF+5J409DIV0O8MT/+hD270DbdgxANNdijwkOsBZOcHj6K6
dO8AINPIsNLIoP0AN0fNI9ZeI4+E9OMhTg3OA49B82Wn+SnUVmyUvpPmm4TrKoZB4DXAwNu78kFO
o+ElyIaa8bJYew2AjsuIFJzoBn1bchjQRUcxK77fVSlpSwlElzGY8Xoa4QIQRsBjnp1UrdPAuw3/
QBA7H19Lyc+WAyx81VhoCUL/9EFpB0xXT6xTBZ+B5nZxNVmIUcF76xqqYBDFvf3SmWj5CBUx145i
hnMPjbHZVtIlOBfU6Y62PtdSpkF3gkDpZqyE4FWY4r4L+7sBPHWgBLZYdfDeyp9K8jtUHhx/Rngf
fwWVSjzJJtNtnqYQxxqa/PziuE7Vvm588w55na0gUz/nCvkuI+7sA79Qb0a4C95H94jchEaSHAEY
FvpsnrFnTWLbF83pmPJTcmSzRmpgauvItFy7n0J26sqPzGBJmU6rkDV3JhIuSr/pGc0KdyXRhshC
1FfAI3WkQyHAKKSw3Ncn5Fvshxa9VAnjWFW2FF4Hfw7LDwhqUx21VS4iPNnPjhED2HOzjWX6OikV
9DJiJySBkaMBdn+lcukk5YVs79R5GVqZTjTWLaD+FDm8UXqngS9XLfIJI+Wru+TeS20mUWbyiD1P
v5PT7nsxCWB7dpQN8UoRFzs8uEPA8hXaIsHSSzZ1h/o4xhJpZVS+HVpHAVcZyW/NgYRXJsuOhG0M
o7ye+XVlU3qCbdwqXHTcY6bzU+R4vpPuLiAiUso9kKN6RqynADWeXA75iL/U+MmsOT8Z1um1I/GF
ECMqv5w0EpttTKWH7UWaXv06BLRYYrmtaV3ljDGDCTXNangPr1Uoh6DdJHdU2+Ns8upWQNg6pXnq
1618iXyIHGTySIWs12zHUfpVb0mj7KHkYN3JZomTDHeaAR4eKvMeGBnaI9E5QtTNofeD/4TWMdYk
NjKiKeleCLjkbIdeFums4hxU3bNR1HwABHdbTIQ3NG4zLWqAjw50uIn3h2/cUTDasrFHVfbc644c
wbDQUOHYxaeUcDBepjyRwA7Qoixg5YVkFcO7GKChAgp/YgM3Wfa+PzuyAnrgQdpSuxzVEUwl6mFW
H685oKZpxsXBIFH7INq4I0RT1TfzzSQmPkXb6lVcw+Z6YNw1kdo0HXqs+qe6UVtI02KzRWCnYxlj
iVAuV3k8ZGQIoEajQZ6SMfYvKCshGnqkH/AW6d2yEphEetQ7KCPng9Oc5U7LZyq1LD+SKGNZPv4e
/83D3q/FyTif79dOdyYPXRPffNLfK2cCcZhCI6gs/60eer/XFz8VdUot6UiKCY/8xt/qW2ggcRkc
QCB2bpJ50rZoqhJ3bSKiry/iLB0IWHnUOiF/29wUFyqEyFdG+tjuZzI0EHOAPeeSVUeDhU0TrBE2
ZsU6I2tL6/nNwn5EvBwivaXaya9kSUTzoCSrv79CB01/9OfejCEBl5+NSPt3zFyDwafy8QBFk/pa
73pwAs9zL/yWiAZr95kmW6MN1MktMJ6b/k1cT3Wm9X/mup/IfVILTNVyxmPHE3Pemm945iRmW2zr
JLURV7HjqslCEkThcHzFe+oEiUccV9tQnShW2muRL34mN0aRkm1Qf2AGCEHlh7FrLtq2RVm/71IR
OXVs64sFr57C4gKsvtMmMB1msVb+WbDENkpGMmgsQGrmcsCM39UB8hlJKcIOINQMdIuIB6Ww11Ft
ynC61ghjg074xxArFKldqgFm0d1OKv6fl0qiHbTnFLxmByhM9ocmS+zjWP+Z38hmH8ozx4sz1g1u
40PFb/AHWVSgy+q2spUCFofBv7z3i9iswdJ0S3WiZ5y30laMSECw+3LyPDKe6mfeiQbwHCrRcOiY
JNIjMUPIKJBYhF209en65B9C3521MnsrZJURl76hL0uq9g0a0j599/xh3ZGee29i8w38bTZXQYfc
XHaw7x2ZwbISAuttiJLMWjpPAWi0iH6NDM3AEiws+NW9pLmV4vMP1FUQmZKTh4C8g3qqX4sGPGDP
sbylFb6wC7OxR8MzBYxUKNbZwKWqyDQ/fv22GZzSKTgDuTV1zkslXnxAdjfoFIcVYhypmGeDl76W
ygPqv/xtze5DnDbJmmtxoSYGQQqJ+BGfELuocou7oU7+UVid3vSkEl7zNHk2ceqni2MnehF4Oe98
qxMwt+x4/hN+pixfG8v8NOB8quiQ2L3SZ4aU/UvyLC32vo2qpjCwZnrX60UAhZmHaGjJU3QWolaE
lD3gwomEc+kK43ZD5tTV+dkt60mhthsxHMYxjMR1SQ3b18BSI3Ecs6BNZllqX30R1CIF5PocAmoc
86EL40k1D/HU4co5zkigNcIqg13HLhBAItBhx3FwzAXnly9Nlfs2CCrRrEwDZW7q9Lu7H6if8YWs
JexrJ+/TebZ5DLoO50XkS1HYGBPpUHckfuvyzE83rlv8gtu+3wQWqG1iJjl02ajPsxRJVxr61W0K
bn9W72XPQv3RJwNAALtjyzQ2t3cQqGcSSlU09JUX0uMSnLQHa9Mr7WSwU9CNy8sfL+mjAb0J1BPu
xU6+E20j76S7VZlQpgW3CaXtNiAieuxuTnWuWMee7TKA5tBkOg7SYHRM+TcierQ0M7Id9swsupEJ
hSG4gs93c3eXPHDqKmMKB457GuONaXK8k/vp4CiuSU2FN81DfvhYnQPBWo9JuQuL34eDRbeJVI5a
5DSpyfqgOw8A2oYwt84x9aHie2ex0SgTCBxmhH6pqop6o5sMeCyQl2oVbc0OmwU2VIBkW/Y8c5CN
YvrY+UcH9XfczDoIYD6Udohk4NXbX/w8c4AY2cxEMiHziNiT7c4+o8mtsg+Ubl8yZK8KOATtfcij
mK7DbGw+W07DSgOYn+xqbppG+bUOW8dK2lBsCs4pzl3msmc13zL0AfR9wcE1CoddD5bFBZdltbo6
K/MqgyX1adG+A4CEFWQPTLQ1dhVWslC08FczgbSGN86y1DHkRxm6FeW1Hq1pYfh348liVBTyLkku
Yo1HeRZEgY+5yZUC6Lv/b8G/gSE4aHS+V93mTtOPiL3sDF7qzA1AyFXwboy6DlHcwblXCX5wQ/Bq
y9clODMo7nOzNtA7k3ebVEf0HhemUpqRXc5K+pTamWpcsrmD/8kn02BamhKJjOgmA2ScycOadMJa
W7qKQKE5o26ZLh6n8Q/hHTglW3+Axmz9aBQVMtZ7vBa9uaSmWk2AJTibxVsR8laj4imz1kB+lHhc
E4KmWuw1z1bn1EFp1DhcIXVz1KlKR+8HHt+fBaSO0u521VytLWtREc5QlmqhCT7wtGvM0mgmbKg5
UHR5q1mFRR31gEDoNfDUpkg44WJN0ZVQu22Rh6XTKOW/2Wix/dhwI65Gb045pWmAlpuqiK8QTo2A
BzIue2CdHh8uH7By5FzevHVH2GePK7KhjX3u+9AjmMoUkPFQi0+QpmFTOqdGGvWlUwwuJghhcvJG
fleHGI2yo1aepJXp1fUzmpAsjJ5+d4g4sae1FVpvSEPC1cMpXqEHyM87ihww0fmasqCDcY0H9r/y
fL4IfHBSdHj77HfJ8j/4S11Kz9theonWlMXWpCYyG6iKgmkzysjaRmcUR1J9fRTqKlTpnSFcuRnZ
DVqZp1lRwLMXe9luHZqgjvbDdW8eoCMkVLBCPUJoJHBhdtSCvKhULl8EGqrbLssBZb34lIq7qrgO
SgQAKlZDz8oKkr77lEOyGEECXzOpcc1UbcB93hVOlO/8IEN51hBlAvjW91ITFcsVoPz1V8b/dQ+J
Nm+Lpjt7+g/Bu8tAKAc/lsJpRcD7mJeFo7i6nUaXQ/l6KAlmq23h5XBcnIPszyYCrFEbj0p14FGU
GeHdWZGI5epH2zX6NoJ0sMmAAcqD1jfBFF+A02UupqhIoM/FqrCzKpM3D32JOYGexWC8Zk/PEzeG
8zRzEGvD8BihDt95mP0bD7/FmMdYDHQQ+KXkm5AxZah5r9PM0Xk9BzQMamy+C72j0IbmnbhM7ILN
GTuFcMNJ+5YFrGk/7Xm1lhdngvpFV2jP43C3mOlNSqkRH4rrkvxPskcgZTVCcsr8VhfeNkcSkxQa
qaYJR+2eszEXT/WV8+7sXhkxMQbIrzw0hRb0Ipn6YQ+3fJoQGUCaaEA9lx2HywRP3zfHOh+dU4cY
BSjyCfaWWkZea2J8BeZ3jiSpNVnpmpbD2EEFisAbunph2vqGHX1zyX/772uLIB9WfGi3ChfU0kpK
yq6IaBnA1KooYuKqYyNpZG9cvTxU+BPsFeIeOSbXJFvFFBHRnCJupqQRoqmbQGkpNZVO7JkH28Dr
FUtMayt+ZTZtcc1EJhyMHu0VaBf7AhwsL68RNZO8nSVYTfin7FP96qh8/oymh5sjrw9UYjAKFB/j
R6X9pjyc3+oGAyEngtPMwpeTqk0SI7aio2D1NxKna7LlR5A4ksOC4Hy19uOZF5Evxu/WXwZGWmcY
TpiRCxud/rcUjuyUU80kRNlkJNbdApPZpXCeGok1FIwBIsdwsJyzpVoqZ22KXKdTw6ShU//5vytg
F9Mhba4sz2nfjgsxOIUKgpZC/GCiDd9sX+X+SXRqxj1Bv0LkSogY1jyMue/MNA1K4vWwGrVV8+3V
PqKeTPCXDFOJXYPB69EA6ddG1NeZD9LdIVwj4kkI7yI4D+pMaUZFUg4CXINU/I9X5Wt0NXdvsSr7
oXLjfVDTSn1B/ZvtP3L8XKMTjSUrUk0MQNSF1GnouQoSeYvZthfbvVffKT7enRYPgqZ1NzpWpdS7
tb1s5hR/juLAZsqbtR3z/tA5xJV+lgaS6Ao9uygN9lhCY8X6Ch8Ad8VL7UpXXq1dwUMYxY46fgy3
bsGVpyOG9eyRuTey+AP8e3mH3xQ2T3BEZ9rnE0rpTDY5m5eHyuW1WRXCJKiZKMJK/nrE/Z1eF0tr
zFaJ8Q7Y7J7PKd5TAzcPG23n3GA757h1MFphMAQzZ45qVPniAiOg9UNPnSTSKuIxHUopbHQbnT2x
dwCJ98n5jHDD+KQRzNeiEFwisKXpcH+m7KDbnss4l3UMV+dVhWiWpGI/EmsvI3JXD0jlyZMJWOXC
vGbV/g1e87Xn5kHnLKz2+tpuipYGmh9M03RsNIU3MFQQweXtYGW3/dk9yYAnhmvixmQEdZ5puxOx
5o8hoqZb+Jud6CTH28dvGYzm56T+ykOkqdz+lh4MyF2T3UuAAobJTWGze7diGVJbgJC8cwYgRhta
Dk//W/uNuwLblTkHhZW51fq+B0+Jk6hiC5AroRx79mn6utRjyZbwwNPzhSidNn1PhxsRL5Twid99
OrbvcXIjnshYRgN40dSktz6rc2B21zpM4L6jQM6bj5o9+pMN2GLjLdnmp47v4gQobPr5S54OBO3f
m8pL0MKARKoL/Mv07Zu772KpPmcaWbnLFPXhK4kEjdF1//lf5hDIDpJQTyYJuqL0Oax228f5Q4SE
igv3L5x27I0q+N7lcwnOIO8SKBn0BFnVg42T2gvQGuDcPwueP2514zZqOPF0Ev4os6FFTuF9XU/7
8Ek0xSYyNEQuDTpKBRXaxRjpNmUw/1StZBhoEmnf4rdNAay5q1lh9wiNg46IKbhHfw/6L9wuvS4g
K1XVSAly8dPwoznCznyQkfqb8X0EI1J27Wlx8Hz2RWsx8hGXXG1LFNGJYVnjmULqdg4gafi55eL/
Oh3/+0eRWPuZvGMe6FutGpx6RJ/xqRUxJ8xhdHWNWUjF3giuYQRsQONVkkEbWw52pYn6eodtbuHs
YUL8hVTUKJIzGL5gmUo9b8kWWVhZCG8gWrfIBLpLVMaKsx2ql+lW9aw/KBGSW1EJgrCCA6OJeZcF
z9BfekZk+FThtNgG0HVBYjOfjYQCw2fynCNIsv2X3zCcvqMCH8MQf6pFYcR0fLjCcFbZbyDHMQnK
mGf7KOJBsauJHMBEqZzSbckZH/BN5WN6RWNfSi6hPN/ElTdN+aAkoIOkh95Adl2CQspHSISYzc0D
zhO8FaYA0IOG8aC111b9SX2yKHzC39cSPIJmmxgNU/dJYWwoSlmFdZ8qctZOyiCYW3CNUrRd8tXR
3s4uLAClZyHbUNYDQR0uq39Sj2efIk+MAhFyRO04ue8lw6ViWwZBUeHLYKVjwuVjwLM/jjnVEUSL
XPSN0DLRn+mF7EMVgrAx+a67wKg3oEkb2tJy11SVv/n6IbUzSKjbO0H9m/6Tlxq7oUAqyBIP2Biq
SSb0Wwl2e3AWcekzN4Z/RPGHB8mNNZLPNiLwibNh6lyIcDpXvb7dd6CUT4FAAOAwioLTlVCh/bXk
eBguNdNFV1jE/5hoGG7WuqMojiHN4YIJ8xEFqO/7tQDG0U1mkd3JN7+TuxD1DCa28R0NEEodQ/B0
X4KwNAtRjAQCUzXM7KIhMMITZYsabVLnaw/g4k4ROpums+nckCr2vA81z83KXLysiXxSE90BWsr5
ryMsWeBzg5V9YLXJcs2r7CxQcQQKv0fK/G9cId0hLPLorsTe2dQ0e4G0jQLjbIgWI4C7VaniaG7h
h2ztyg21dWrz5sxX4Q04Oid5opiZ8+Ft6QTJFFkgURmV8BjVonCXfNSuWSssRHw5z4jl6g81Utvz
yKDTtgFW6CxW9y/Yf7CxCYPfiYtqUwGvydsjP16zob0gUKq4++t/5XLvFHPq6Fl13DwQ7RMmGwb1
3g4ApKx4E/rkaBo2kYbU83ymLcqJ/NCES5OW/7inJ2ArJ9lXrIG4slK7dPv9LhQ4v3LA610Itrda
TDWHfm8tM55xXJGMeJHZJtfWuZjkn8ocHUy+AWPhAhKnP0NuCEzLiGhjqPiGKuPYbShWOZ7jiWiD
eTmL/gP8SdA4bihTGmAOGkn4B8Bmxl27f5qDx6TDwKd5xM6nEtdyNq2EFE+oE1jmW4ZrLqrSF+9g
GEEwxOegnBEcMUSTtfevu1cz2CJH1ioPoMb2kvzZ4Mq5dOzPS7j+7FXA8La9O5W2ddCEk9sLJw0U
b/kTGlWSUTZmmwXxfD3HZiws6kthRPjkDAUtvSdcq5bBj4276RQI9gu9pss5rm0WYTrzvPvcMK+k
KYri3aUNWQEgDwDo7427USUv88vNhgFGg7MhXXY+5YwkTlmmHyRHUX8E8go2eRR3DVt8j5+yeaJV
jq/zj/x/GZs6P6NxUokoB+Y4vM2asa5GJ3udAXNz+YMz4BjCBxaerzHMnrl8mN4QVV5BrZ1M8fW2
RYCxekUGZIT+0Dh+s3rCzeyxgPXZJdmY3VVwx1sIB7OjTdAFTbtoKSZfl1u1iPb2zDwU/SUbKI6A
bLFZK0vJfFegtuJDqjs7zIPyfBaDVNRcWat2bCg4eq24Jw5Mcb9qyhRESVXtKYX4JVQDhg3w/uA4
V/ltKlPSLjhleCxquOq68BXfrY+oqhGt3zCcmsImtnran7cBaY9IOpfkobQkZroKZx1BFjo1cIln
g/9QCulD1XJY0EIJwIXhddrB26/NioOb2FxLSq4LA8AqroU0LcaVDt9mP3aPRWob1gs8WozTunYx
Ihx5GAhB7eR7drYe97e3Pq1oSsX+dj/uHoPhcwdrsftuzER1GODfwaMQlE/O1J1yg6tYAhuuEEOA
m8Cu7NBQOvd9XcLSASG1bjjY2rzrrTHYJt2dXgFbl2uUunVk14JQjgBh7g5KiTj42rFENsuLJasw
HPv5sv5DtsQHMAapWmj9xVTbHt6E/JavMNVTAXjU2Twm2SHkDrLKSd+5+DWo0RIW7e/9G3yXsvVC
7T3wjSUVZkt3xp+aDAuifTGTt5VRfkUwmlwwUncHDvEevygPqAn2t87dToSqKrYBXySVl4dqU2d3
FU9+KeaP7vHEB+77u7t+JgrzI7LnaCavmtOzODl+aMT8FaASy1o8PHxF+jBYVrr6rLSmOf4635+p
S35f1K98HGCSQ0QTZcQFOPweJu5UScl/eRA/9L5R5LliFr2uNNYm8SSwh+NqvGPTonY1Xw2rpDpm
D4KCH3DM0/hxVCLU9JzNIRDosMm5D9Dn9JcYewvzK0IJqXqp8tbL8vfCa4tyobAYhpq9XN3umhGR
zMJf6jGUtS3WCe3/rQkw8D3rB6YZLiL18XAs9i8gUIJUHxkYpLdv73VWc3bdXA6JPcntiGDUNEDW
8rQOjQAQ6FkafEWsOhxCGPkDEem4oWgrmefWRScUmi1s5pcaxfNfBakr26Iy4OWF2SBMAj29xYdH
waRzgn+l7NwKEtufg5c5VrnengSSVC4xDu4LXhS2ERRft0XWDbyR4BaTurqtyeXOqWsL7+r1dK7H
JmnOsOxmnN8sz8FlBoTu7A4yFQAVBqEHTLB3slwjh8sv5+WqYi4emuAgcLzubCyY9kRnnF2BvcCP
oWnmc/DjTq+WRfzdik4SFrCYQDtg2Al8xtQOnwV6noO0Hp++RzAWLsX7TVeK5QQemtjFvagy3dMS
6W0aQfPjQfwHoTt1FO1ada57EE3WlvfaMEnIeBHzHCitNYMj9jbHfqOifut77x06xlmza/qYFWvM
ZuDCwsDP2hbWAceYUvhV3xxlu1ITeYzYs1HyLAUZQj5H9jw7wdnlKDOwvn3qqz3m0NQry13dVqM1
QmOF5edTKyvYp/SdqlULFT8AIlK0N5VXP2vL94A6saLhdTYno58nVsOTCSxekLVq8rhL5t24rbI+
ew1XsduJbw37JvZ87w6bAaqp/EhEx+iTUAw8KlNroApgnHxPKXkGqI2gX5RYB/oMMv3poA17UNob
MTC6+Kz1DUK75f3qkkLtVIZlECPy3g+vTl0Ms8mP2SResIYboWy5xCbVMzCZDoUxkmsr+HL2VI42
lpUCU3g7jb3PBbcULwJB0xDewEFAL81v1Sb2fOCo7L8x7ZG+r6axmcl4GEpZbRjOrhepP6ztTdGJ
XhRcafJ6EGdV1aM6ojC9K5w7LRhEodpagWXN4AskU9DXkZeqsAjQO0wz8Fv6FPF2BF87pT2ch0II
wpXfKUgZRRkmLCDuFpKlDjlfHS+YW8ZYEd3m3jm+B4c/b4GlQFM15oGYBr12VP62wYHr/hr3A+JG
GiKzdTj5oOQQGBOFusE7ILnTCOSIEGKNlS1ol6gbJE8h7ymBX9Er9Z/uk6j+3fpoKvph85U81VXA
TBPHLOksWXSocVZg10/z4zwOli+woBt/vtS4hkfAlPu0aAJw4JcDj5/sHMlHGfHTvcCwUEUdGHke
EqEVW2gFIIIwTjnYpTfjvGD8XyWZ13AjLD9Hr1jcbxWRqTW7DMbpSGN/gWHsMA7gVeXANCm8pWna
8iWKONAFnKFcOJPzOXfEQlOseIftSoeTFRHrHcC/81FpkpbVloMMF6x9AVLjddGHqTvJYdHlDQ2l
6JCiSOGDfNWz7FJL0uQP3Rn5nZw70Z7AnUcr0Ym6eqWIJQx1OCeaSsKvIrwWzPhPGVyk85PWGX31
xODvJYS7ZbcOZIn+RDBitE58BDFGXUYWWqIH1Oh1O5Em7obP3gCNKwMmJ8CjhsGrCkqIsraYPCcR
CEOBwry7vwdh/dxoDQYBEEEH/rhXFbfTwfYnruoRqoonUKSyIgiQpV09E+C3d0BZv+4GU574NcIA
icatERwBQkLLcXfI9SAGsdnFiEr6XXZyj/+Gp0lNy1pQjuBC5R6OUZVAfwT5ohaomYSgMVjWa1L+
p0kZrAQxO1ekc1yX6LX8ix1MJ6XUdJ+M4UUyMm4+j1UtSx+M3Cyk/vQA+l7C8bB8W/+dRFjFMip/
LggUbeBOwcuS7/KyZSSYHA7LSu1ikKqtIzcPyVNGC21WOyveKNyJiTbNJAuUFYTKFVrM5RTwR1bz
dZSCFi/X493+50E0gPc5YViZPs89nVa1Y8Tlo2/OiZx/c5JR/aIQnSmfw95f+ne9PW3+mbMe8WWa
1LnED0YRTo+DcT1fAJpMeovb29wHI37MvVSaq8Esnc2PpF2/qndC2mi+87mYaFhAn1WQVmG5Xa+C
fgN4aLisSkVuTfIXSMiM3mmVcMN9tu/1OKF7ElQ0PAZA7tKrsZ8kWOqPE/Wz+QAlXPqAYGb07gAa
+RGas/HLu2ciluumT93ykdCPIwD1FStP2DThwvOIFv4BP6S5u2GL8jwxsb0dNTNUESgkKgSA66Vu
n4fTepe+Xn39Qm6RXQETiHbYTQClyJ53pqoCV9ZcqksNtmF77n3sprGi80Q73YTGbVx7djSyiwGy
r9ujx7BvQjSY3FH4wq5GYH3+n0TJCgVaNpDEKM51/G4ttnGBcWmY9NIVTn9loFT7OrkKT/2Deba4
8kd91vuxzHcy9bKtROxbPJuHBmdf9BMlANESg+/6niKn0M3xOoz3v5bo/GZWSFqOUMQUaJn12IAE
OMdIWtngd9Wp/0ACzwYpteQAyjis3PA8gkG/t/4IRkl5KuC0j4xvSMn1E/iRD+gHrfvrpUbUGRLK
h7UL4124NEF6gTgOa0l4Pd3TM0jTEQqi+U0N6QIBwq2fEnwi82Ucl+cn66pwyNxvpwXxSyQmmPA9
YYbHsOK78SZpIgUPMW1gPAgj4/68k3oef6VvUqHv03hsXjBc8enkHPc8V99pQPjTn6Kg3w7h8JpV
3EE34bPR2U7oMw3fv1AFVFDPmC8aFke2QE4muVD+ua1B+1fwiO581uE+wLnA2exFHcnMH0D3CBkw
FIOkgRdHHJT1U8KUtqs/teKR7a7D7CC75S9cZ1NdLuUsoyJM/SMxTxDNPUm4FKmCqT32Ia2LqNgv
gbIx13b7DbKOSDvJeKCzfcmkXwwbYPFc7kJ3DWNAxfOvgKSHLIqnSkM91Dyj6IzIO2FmTjGC8A4F
WewFt478Y6CUvnOIBmJwRl30ReYC7IOse+xj5S7k4GsUDB2F1Np2BcYfgwTCWBN29722YjVGgx22
c2I16Xv1uci/TV8JCk0ocE7V0AYMnaJ4B5gacuhrAyHvnp8Q2Ci4JOciIF057sJA+tAuXZpW+Glx
QcHd61kwGnK10/ge4xntzgouO2ck344Q9C1jvKfNPnH6a3X7eCZ1RPPEkGRZfr2v2CTvjsEzrD+2
011e+HQHzD7ZcqP6/XVvNqAYM/piktG4ykUqUu8Ff+UiMr7R6OodHdX8UPJ/fPpc7PTgzzXGk/o+
iUrLB50cSk4m7KUMxD9Yvk60legB7Xh2ScX55+5DClIcklpVw8RO+N1x0YRnh97bn/NP0tznwdBf
+9HkFAtg2kMuEMdjGAXnC4Tl2t1TmkJ1BV3kuIwJwc0eolTuOmgJz0ywnv46j38dpYIazsvEPhch
QzooOXlloQxslIqhZ7ZmRmkpiuUui4zHnEpuh6uRbrCT4OfDc2CiRVNfbUz9sLZC/9TykgCH4rbZ
o2iWlgg7pgYv7AWA7FSG5fYpoQPCmEUKepRgiAZhvK7uVk7hnfdo3BMGJaUUyLVlI5niY3Bmvjjh
vtorYF6MaAsFCyJE6dNIlm9jfiqSHEXdKDeo2J1egI/bgt7mhaYdLFMeL4XJCev1GzNv83vxhkA/
/Jla172Juhd2YoB7I+m7y12Vjrf/cUoY5B7mlWkHQV5GMHaKY84FBiz0j41ljeVSVdNW9o+qswa+
y3l7Yp9eLoQFbheIK136O0Jyh+qlvfUs/cGy+kzBQsSTFCKEBfBScH7XLCdYuRkoK3L9KIt2KpNj
D82A/5hbQumIfxNsdp2QEAxa/p0fvXgEgpl/6zR8VBgmed0CrT14CczIUiOYSKnhkx4SCRM39Yu9
TB43sMqV+CHg99OQWySHi/TaBpY0WXtzVRbSbH3aoauep9KXShpyk8Jm+35F+/aOiOgipPyydZL3
NSyEoqTChXoTi/E7DL/tsPOpAEtaqkuYP1UCxr9nyax+Uy3+EmDpyocTUBrQHwzjc5UWBHyHDfsE
wLBRisuEp+FOZW8hR4V1RACiSGYXhR6XlHT0m9fQ/HNnw+NeCv9pKKVq75nd3YNT6JVzfAm5HzuV
M+v7DHHSHbZNK0ui2IJFyet8qgthQaqxQNwG7X9T7RG/L+WuFZmdBDlRjUgCidpZq/kndDvEdI5o
P/lQbssAgrDJY2bby0lgcE/KVxcKXueRMeG094HbFsPwGtZ/5N8hCrv/WfJAkkNbLzPyh+/1x1wm
Ttfrii7ruOKkqcAZZQpW1y8WTs6q7DImMM00qytGbDM8abRa4XbOhBD+9xbaZARUjOzxyd8nBsJu
SoiEVVh6mgQMlrpUWYvfKI4ZhsGnAmy4chESYgAzv/CVXoNvVSFCpHc3IPSe29PxclxOk2sNwCaN
8O8MhbXeI2Ek9KVpSPLsylv/nJ1wvWVQWJDnZzoJKOUt3fsaULza9+e8wn+YdfWKwXiKLNT1XBOS
AuMJiB2JdxedU+7WiF2DGSesaVmtrxTZagaI71QDGn1+H3fCOYg3NLnSB7Q9UgOyiE6sZemf9YOu
S79eC2r57ldEnvVCah+T1bunRJlfHeIBFyXK3K+Dn+U9mgBKFjWMbps3leKopo2zi00hJI5TEGOo
E6pNAoth1cn0GX/xPZ8ALC8mKsJZuImZ2ygBcHjXe1MfD/9nL3chpJsYxfHWrZFbVhMkY/UWDBW1
kUPW23L5b9qUq84iVdcwegMzL8kmuMD5ip9o2a/ArdZlVy511uhznY8Zz+gd9j7Z/XTsMB71gtdz
PsAz41C2JOW7KAbMI6Zasyi3F5BLvcKH45vVUzux5IEP1lI1+rTO770BYtOTfUk7GhvOr9OdAYcf
rEoA3o+4dFi5bJATDxt/kTaV4VJcWKZ26o6rQfprPHFBSXMmryU/m/53eXyUB77+XLnPfzgMee+I
9Wi8yumG2JqR1t7AY0eCUuwebVES+SfZZYG+xUfAnDFPkp6yFCC8XWF1iQrwWy2MZYvW4ZfkAbH5
1vdS6U014wHfUJbtY5VmaL9PdZwM33npsLjsGF44f97aXDaUMPJPBLB1Nl9oxCMdIzagwkS48tXq
xRRmVybvTHLmkB6rUvWWMSXXxGgjql0ooHqnHowdIYk+sI0LAF0FU+x4yZNIpaBGRquW6OaAnhVf
z9TzpCkYv7/Y/q2xbF3Ec6jqOZt6/I7iZm8lWDuBVVBgv2o8BaE4sTYRblJwpuv8/V+Jhwc2Q8/E
Ua+Jtav+esIsud9VgH2Xr0xQLzwjRsI0GEn5wil3SidOht9XcGJTzIWkaAWT2SPt8dcP+ogdfCpH
65CLXidz0Jfm/W2hRvKcxdCa6LXkGmhbwtXvlhTxptzxIZ3uqWddW9OuyxTAWccmw23OePjFfVcy
dO/5S6maKz0BEtS6M/vPoHxwZAwd4RmmF1BnCmAPtk6wpvATB7qacQrDHWrr6AONkRoUGqQE+EIl
3H25k7D+FaZMNkvpFNB0JOmt0D83ischkUqTFnK0XHij8VeW2PvqB16A9wZHeMqUYplf1G3HpBrQ
OMJIwZya2a40muZaVLiBaPSMcK6BgzUMR8YFgPvHR8V5A471Ewn6qwIukJ5XfmyT9OmL9l6G2e4B
hgIKzweACTStW3aez+amMt13Sdiv0gAs2bwBup/fQAR7hDnPpdJypn4jTFrlwmdVNsY+V0c3BQJa
D8hFkOIX47C6NCz5uPhqehEt1nrp6C176qzzBWpPDC3bZZ8hBeiJ74FY6sf99Hu9FgLQWjGPBZCR
aor8X6gxKthJg5o7/k3JlNc8fmKrf/4oevi2INYpPW96OghWRhJft7Lfuov5GMEypCJPRc+MFF/n
QW5fsi6BqyI+C0PKdzQHbLGaJJD2UNbsLcOj7Z6WJeTqRDyUN+ynwgPdofxMNoXp0W9yww9h4Se6
mGHUhZTl/hdbNveqsSdet8Ct1rwZzNOpLEackag58z+wwkz5wT6WU8YfgVyAAUlyzFawV+2qJj+r
/QyiUkxZLinEdYZV8tJdqLxSDEtNrFn6+w17+qyVc1aK8NLKZnRei3gVyVXzK8epqETiy71S+Tnn
qgS1ALJdYvET53IGt4DCR+xx1HBk5Mohiw+BLfEHWY98QJRMJBah6LcEb1eXJqGuqyrl0BjBriex
RIO6cjymR32NyV6OKRjGm5znvuVL8/tprDVlqq3BtgHzEEDMxVekwEovvspXdEr+h0nxceJjfevG
6lJqwQWF/3Scf6TX92ZL8q80GTMngk14tI3MG6YPlbW0lLxZhyQllB090dreS+Tj89J+TBTJMuOd
UwmH+EsA1X77F3S9HyCmJbTFcHX8gVl09fLBB4Go5Jmin4o5u/YfSWmrzjKoKeF1oIdtcakcbcme
i6D0BhTpYsI17mu07dtSuKpmgXgFyhI87HO71lYlCQSTaAHs1V+GnCheDpM1TBftwyAqL8gwuZVq
n52ylHf8sBVoj5AgZ7AWQppJOn0dCHrxSwMIes4uiWKNFSiadS9AOMf0MGsXgpJSZvC365+P3Ujr
oFeawZw0j/yb9DHHOg5mkRMY/7T0RLRoT93D6blQPNqoTVHUQdwwM4juuD9KpNNgN7gt+sT+izyt
no3DHbK0BH+xyNWX2f4j2UVvrRyBEfO4q9m4cTz+w6NfVcuBf8bZD7ly6HNbor/Z97PUURgZQObj
gxlDPVeBZPeWQwAy8zl+D+uSgua8Y7ZG1KrhqbqkHO6Ya61C0/5ELgDnqZ3HwWDZQJJKUqRrU1oK
0SD3hRXALTKueIwXCYwEwL/rk0pFGhhlWjzfNMHzqV3Kizze8Yw3JWq8CYGONq8VOaxd8FnAsRcb
EW3yyGsYGHHdHqQ7TYDIB53e911c1wihksR2pDCvKP4R1CdfBlL/8eUj4BJyRi/oGk3I9FtzzXZX
jxdKnb5u+U/nVYrPEoHuGQEUUVwkhpQM4wCzOUD/johf9wHQIQ9uWgj+za48IdhVuYj1ZDcclioV
3alFoVtCvkR1e4xr5gjTMZNfcmR/QOyu7aLr9rYn3BIPxA/70eLZBkGMDNpgGDv2FpYgtklSsR5E
CaS1cxTxDN9Vp1HXxGMpTunhYMRNZcTUxiAa8IVuEEvSb34xqVZZYPu9LtyIK6AYXra1D08wIk1I
FBqFdfv1zoRpqsAY/e2gqTzNvir1j8KPOEcwY2ltyDe3VW3s9VcpZD4Ml+aHkAL1oN2lyv1oMsmH
22gs5iFwn1P47LEtNnTgVIek/UMGPccheTHJ3Hj+a7CK4BMcYX/XNbtXOpnulS/u6VRWfTwvOC8L
kXOvzafc999OOZDj10ZPYeLE2dK/fsh6TcPaw5ZbKfn8aTTuZGwmY4HzDpuW3XNg00VszoDqBb2K
4wOGmaTqDkAypzhLYE7PJh173cjjnbr74YmhzfmOs9PycQYXLNT5KIoOIh5Qal0+6OzvB6n8zjCU
fiNTwmom2Mr4+0YSXJH84nPF+NF6D0IbySSrnXzFwXfUZPJmwWKC6I3ZFcAlRJzjHA/lXQN9L5ia
+pRu3Q56xRhLl0gwljCARz+EwViLBoGSBFVkpGwuU9xih2qtXIxLULETuE2DmB/9fouzDCYa2aA+
/2onf//NBpZNsb8uzlYmkr7Hax8uobVacilmO/1yzBWfwgMJaAsm+vPgky1sAp8cWe4eRk5FxpOp
kNBCjp314zZU5LJ69xU5WnOtc97SHmNBbILPtilLOtoTIKmlhyEeGmNJvAgwEyUok5Adh31457pZ
fz+8N32S2Gsay7XqYoLTEvHClNwRb3MuUIx1QVWNPzBVT7EXJbb5Jip34lN1r/lzd/ThHGW0X/z/
Nj/MOusNqCb/JDpYmbomQpFpByvQsFxZj6EStajk4/QpUZr0j9/9onT7vgFq16b0811BuQA9tRxK
gyXsLLN8OOCkPYJdCIvEEeclz4zXbPKfi1uazkCKxTzkff7AAof5hHfQmoZe/upFGWmDxzzcfZ2Y
CFE9eiFBFo+7tCx4L/OLrNd4vLbkcrsLWZ0UJnKHOXliUS4TAOAtFmdQDvDejE1E5K0KVcuLPrYp
CN3MHNih349JTYxXkbt3ONZsg5LBtT3KmCTnHistl3ZK0s9kdlp55cZV3LrlEN9t6PYBbYEznxNF
v0ezpz7KZljNMWAEBAdR8cDUVwPpKKWF6DdaySevK+IlISDzZ2btLgTUXrX2+nt/TxefHMqxfIkk
DlQjwp90KyA2V0P8ZQgZyd59kSBgK/8GHiK9LlYjU/VPcSXTUbfKKuQkupIqie6Peldx3HKfnPKC
H7s4wSyIHy1CJRL9pMLrB9lV2Dg5naAquf8gK6BL8O5e61OYH6SLCEU4YtsX+yo/AkwR/0u8kLEB
loSqtl1Xjmalw5l0CE1447XnBOAy8BsjgsC9uTQy8+hWMeX7btfVxWreclqNtVBjFSII+SNAoFfV
zcUTg6+HHx6MQPwvG5KUCHoznu1tr219aRShOMpflxjs7zYYltWOq9lfbGwnboP3YXnq0TQFaqG3
GhkxrahOSCCLnyIhE0RG6GGspoAxsj14Awt39ljg7XUEPY5oX5Y0iod6Oh4ri6ItnRXdADu64OXC
9uGbyxkfCv73eH0QjyKvnL3/zH7CNFXqyPgmRw1WYWgUD2goYPeRHiliMxaUnxrJXQYL3mg5SCBG
oPlxLhAgM/bBDlJ5wJ1y32RZejwvVQmxaxcyDB8SD99rLA7r1JxWU1gpNMBRUay3dfY+b0ayBBOC
7EyuL6Lx82HDrqec35ELDMXsQbeC3LWAaZvSgf8vHsqISollsw1tEFN0XxIwGXi/flkzR0QoFyX2
cOj3WVEqNnbCU8dzkpxtHcZgpTKxniodlp4MMEcMHsqNYN+IzNY9arI+Hm4N2V7sS0rbGwPFkNp8
42Y73+B7LivMIi7X6ds442zeDn9zMx8K4cxIF+Rhp0VEme+d2Ljsv4qZXMIo9ggYyf2BXJ99ZcU6
tUfD0mcU2wTEp9qofbOf34VX4IO0VGnglebZz/EM1vn+RS1INbzMW4KGeVyU19WLQmD0j4aSy3o2
A0UFVoWKvqzRtPDudln2IeGYsVUYhP+fTHFhYSaMsB1vFIEuSWEbhd//r42nPL5QOSQqwwXADkSc
h97wCKTZ1wp7NkVjAnclqVTsbwXW3GiC2xsUcVszQPiY0tf3zKONp1zWw9ChyzNURk0xMBfBlH/w
VevTBe78JPGaWMxlYBX+HaLiACzyVO/unbu50O9ejGmZ08PXkVaiqKEWG+G6IYz2K4xcsGi894O6
0xp7HDjVotnMdBz+qt2lYqLUpSpgjg4TRv6hxolr22ReFG6+1I3DWRF59ZdZv3C6yZBdTM0aY4xR
/mU1NgBovTyjhrJIueNvEFTEqEW0zZ6zdPvgbnNFj+PoDkXaNMB/c9W/utgsfyLxuvMUNAOCDEmW
Bs4Uaca2loRk2OkQh2MA6v6mMwnhKQm+0b7sDJ24QlqzvGD5i3To78LwUVWieMbRVwNksRJDTJcw
LVb+xRFatb1okfX4wdcFgLW0Y0SzpPl0vJX9xfPtXz+o3WkllCiKtMG7ZEzIikumCnfBVMA2NYds
vdBNPaXPDcKwgoogkaJKGraZw+OUqpC2BzETGpgACy1WnMkQshAJO0LOdlzYu8H2XfVhzysSVpLr
ka4z7Kx8caVDUE3w1Gou2B72TlUzktVo9HhTUAF0TfdFX4SSzSrllVISHDo5YNx4e+VApl6ou4Mb
W96qMenBxduE6izFGGlwTwk3adZ/al8sXehGWzKsYH/90xBTFVeZlTr1x1k5I5uoSUriCy9ro0Of
l9dKca3eJ0OFioqlrld020YQxwFmlj6AIvTtNrl2lJygtG7656lVYTTqhaVNLORSp2dug32PtErc
5hvQrT3VyjnkdKix0kOg8sz7oVsEW9t1G3ABVmQbqgtFKr1SORlVHp5BnaJKW8uOxvY4QxvkpXu9
bQpewT+LSze9zd14kAIzvHBYsEnjEqBMZxbYqR0EsrUfC3JHzB0dfU3DtNmYCreoO1n4BKfe5Una
YWiElxHkFE0wq9wJBlpE+AGZntCqwuon+wO6Kzo/JixV6sb18QAajCk9ewhXdGgdYUyQUxN+rMIo
v6NTRpGvFwnFfTVq6S/ieTcjuyka5Ea3GpYpM2emNamAOztK0IV4D/dv2pq8QB81EbPF/GBZq2V+
zFcA6C1Y3uQ+osnC5Dp0ZlXV79MlXdk44y/GIEkLvFb85YbXoBbYupVYFltdHRGFShPuInPVmRJA
YJ7QqP9b6zxPgMq67R5L38/0Ppo2sytC9EyqYarDxj/ByhaKhX/gt2ZdFMxjvgMqg4Iwg8/e9xeG
RGcNBQYKH3joxRPhF3VEa+aD0shEq2ebuZ+90u7YTkCBlCH2YQ3wS+DENeemgeVPcPMswpIi3glc
MTnrqCInWE0QU5b1/Na1TxjM5Z/WapBIMYMsckj+wfy54ZsXXPGGHRW9xeboOwhOLAUw6aireKsY
YdUYrwr6smugge5Bm/4CBnFStHTu4bMnfALoL2daSJgpQ5WPU009cylRre/panFeagxFAjTZ0DTV
q4Pk9AFF6jDOid+QevU4ZrnJ2tjamvXk/oIyMXzQURj9xCoQCTmWoZDEeWwQBPUhxX8QEO3JMN5g
hf+vdb8Fc2/IAgB3wpP0UusNlwSm57f9BlmxhYInEGa+d8oaBEUnAAuWpylYdJgnVi/BmQxuWriK
UrAgcX6/TxHGb+E65+k3K+lXKG4lVlHRtUMuUyyIPbekuyy3ZoB73iHlDyV9f3Cw13TTy6JEApFs
wEeE2jSD9Ftv9z/4iUatAnUbUv1aL8QBgpShd/7yrcsN3kiygK+e+gzkmTOsAMtc+GjoauaeF+On
BmLogqKot2KvxwBwbrtcdf/qp3OOEHbhq/+qYbSvMHdQ5PIdv1GBPxtX4njcdxfW9SsexAJ5a9tQ
ap3kzcjRn0wxgSpWhNz32iSn3ueihoKjdOvWagkmbbw9lPlHiugPiZvMGAht1o5A6tloQZfpBAND
1s50CDFwOmb4I5VYkqpB7OrQUt0rlBWqvHtpnJ4GMBnaRs3uyqIjBROzfIOo4K3jSa33rvw9X4Dc
U0sa47/wPA2j7gwOmc2kRj1WmN+kms+J0Iw2Zh2yetcmXRSwLaIPrCCdDNAg96kdyC/jfuz03Bhu
V4xNsyBIF/lwi6gQq1IRQR94EDXx3jLxJv3zCQd+BkKDsYO+AasACvjAjLBgVOjpGfwksrIGf9cw
KgeiU0SI1xnXV8U6mTUl1gZVW7q90TnMTgMP8IHnnFhVkgiFgI7VpM28Wachiobu09S6YVFOEc/i
9sTyEQKNFnrPEhZ3kD6NQIzSKFYBgm7QGhI8vNrHmFidttOv4opFA1kPnX43dIPc75WtPiMz6tyv
kBIlQGRqNgiZw3rsDzyGEk7d3r08fC54jaqYkM2zLQ4yuGMLdZzpAU4l8E2HJH1e371Yjc97hdh9
O4uld7I9xYNm7HGYZHeozcuajsytJC3kvHBR0wgw8YCxd3W4VYSnUHRhlA04aD5uwFvIR4Tgvyt6
xRM/t6OB2HcKT/sdgY1t6F0x+Y/oQR2Z3DiNy5XOar8jgbEBJUKuX43STlzdqoof8j85AV0JPKzt
zHDk2+avI+7gN4jshXCwrNDCixjiSTyJa20ENqC2o6/juOJUhGlUGQvHJa2dKt8CItzVi/fLHaU0
bgMCNw1+5UIj/53fn6Lr8OyMT+OvLIFs1kbilm6BXYHHb4NI5z/rOg7unMjrmYxj8H3arzi4g0zg
lD22Ett8g+3rvgWjtIYHVGBUtakLYODbya/n1d6QmVGeRpwaQR8SfF/k2U+8I3++9ZdB3yjNNV7v
c63SEy8nBepYb8swuWS20mHdxgoP/T/dQ7EGt/czqVmvSY6hUFX3lxBJ7CI+R03eEYK3aPb61vKx
0kNFNQVk+rKN1AY9fQwbgpK9MMd8DuhO6cYqDYkf8GXvTv0zQpd/q5IIT66bMkRwShLNzHTMP7aW
Me/8CsJBnIcOM+ogln/OEkMc9waEy8C4TJHGDlgETorw8Gko8a7CKuTwpISE7QncDQB+VmwfUvtZ
MpphcZVqL/jeswVxp+GjjDMMlEfQD5hrGUDTuNy3yQZ1V5Hk5Go1Z1GUk9dh/xgr8tUvo9pJaTBV
HW3WxBYMgO10Fiof9+/LCdSIozwXAgE3oOHGaxgOgH9gKmxW5CZUvc8QAlgyK5wKnG2zZq4NzDjr
BIeukUVxNH5qISVUcR+6ZA429TdqGFC4HuWI8UxXPAnoWeGoA9IP9fkpurzfU49lSGazpUA2rOT3
wrW7ebvoV1EbJ6Tjt4ulimN4vhbhQqVayrdQa8pK7fZfbc8C85cFt+uj7gGOgqy+Oct5Jgn1OmZl
iGv09Sssj4yTqBHByPVTOkAmLvNzd+5nvxOJ1lwdJutF3iHofMCEybazpYrk1CMifN6aTyg54OQx
g3Rh1XlWvtXR86Ku3/M22ddkZyjhsAkMHKuJhU7nKl48P6IDowekcwsy/b0TrTHWffvLReeO8Zkx
cp6Rngw1uW6J7dnIc65iT2nnvjmen/nSCGGrqDweHEbd12pZGnonP/CU27U8m22EXw2FRKDcQD7p
GTBxECcbM4afnbtblK8mRBcvPyXJ3ZetQ/A8MFXy8n/awvm5YFWBcyZUEOI4V+COvVqadxBaXynH
QeOxAzCtYznpPT6GjEn3izf7XtrAYKB6RXALGbfw8URu1e2Ij3XxBLtiau2K0GDOcMlK6qvnKwKu
gPNiedboD2GksUVYMwlYWgByh1dsKhihN/x7mHK4CSQfPkLv/8a7KihYcdiV45Xgqu2Q19gy831m
YLYTUf3ekw6UfRhPBRmOrlil+Rpd3c/xoSVL55cRQQRCIQ4gfyfVcNMkPrHT/34c4nQ/PqnPhY91
kEMGkwCOdPLPFkrEPX0xglDjZhAe363LntBiteZscl+2n6Nlhj3FRjKa2SKFoiKQ7IxAe/TTUMoI
sWZzijdW6lhCbJRyjUDbl8vuximHU9L1u8FagJum8/yvNsD1vttWAB0jvcF+rjqKV5ODj9CT8pmp
oV48QcdOdd9cx2vIlc+2imeisA/HlIn0cD6tP3UOcoGvXCgEEb6mxL3Ia1iDV0sFdQjZLkga8KSE
ihlAjhVtJLPYe5muC7g4N5OG7DI+0plB4CXARr+fxKMUaNveoCAWjMBn6ZJQHJgWq2D4CGup/bcd
t8sasiCQSZkV5+D0mLuTKi0MmaBGbNKCiJ+P9HaC5gFA27xaPKZkP/120GErU7kJ44+yBa5e1HSK
cMCAuOcu7gGzByEhLV0gBHb4BZaUR27HCPZdO2sbFSZna0A8LKeWXgka4RgBzL8bFOIgaqumlrLk
yU/mgHXyriH3MkcXO9q02P9XKy6yt8JYcJStbnusi5c/zKjozhu0tZuMOsBl0Sg6CtG3toKEFW67
+ArCHssasMMhdJ7qEki0Bpt+Xn6JdO1MJPNLz+MJhAI0YL+WXit6Pg3/pbbA2bELoBRQDZ6VL77H
PhnjtBElxxWr+K89TvY8dOvBlQbxr1oBBhR22aQEXtcw8IKtWkTOOhxSgI1WVbkgtoOju6wQUHhw
wfiCQhzGU//4WhivGNBWmkM9TMci0jMuXSfXWF9diFnoEOn5V0BfXytzpymYVhBji9tRsLmJ/k+3
ODhhhHetOHDgIcihl7vSSccJnXadaY+ntPIZpu6AYKTUr+iYs5IlqXe6q1hl01M5ZLkWuEP5jpa6
tDuNjpLA/gLfDvBGyXiPocSaX9WgowNwXxvNXsxXaBrAZFuyaAetQ7FKx9Sv0wuPzC4/khy+ISg3
Q6jzo/m4uEFix3YRA9SN7uvZLxP7jwaCRbQqT++QtfPKVCe/0T+S/Mlgprrp8xG8ldwsMB1pRguC
l92dA3g3KAehsL9PlkeCHNJvoMrMAArdzoygpDeE+ZUZ8Ec2ErGjuQ1i0tlhjAGAl7QQmgeeW19z
5He1KvWMuHAVmJpzgXF/beW4uBF6RCNHUGnnAf5FGjFFvIjgX/wejNC2kWpeV2uftS3FRZUVpmge
lle6nmQHtBGDRsbJV/IwtC45M+2scS7d/WGoK8z3l39goT2BNCi9dUL3nnusuRue7aDIWr73UB0D
eLC8MHiM+f8EqOd8HlGS0E645PqqmWgyuAH6jAX1h2/iXwYfMt0lk4t4aMytv77RjzlDozoPwGhk
NMbVBgbpEwsb0pWy4Lr8S3PVB548slsAW9aNQkzPm3me8Jded9Jsk+EdJ4UPHzCxDf3cpFXf4+k5
ITlCRpc0Lu7Rwaf+Bq4YMJR6vPkSGxgyST85+R80WOQ4w4UJKoT2dfEadkTcseBgAQOFHICwsTxc
xiU3yGXAAnX+V/V2aC9458KRf4uf+kTOClywnZDr9T0Q8OS72LEcaE4qAhETymbCVGll1ThTD3tq
ECMYrMqb99Bp613Z4p4YJ2IC1Q7+W72YkCErqatYA3ZhmCgvJw4eQdrelL60jeuGYlz2yJCxrfWS
lUhFky6VcIKrzuekfwN81L8bfUz59rlZZKkiwV1sJGs+RkUwf2lYLoPY3MOQoC9w1WWlzaOp0krZ
A1QayMYUUjFU0UE3NOWyNskP068Wgxbk948VDAkGMcdOjMqfNjDiWJn4ghQI3/YLIYmUhPXZBLPH
qKxSatAuQkghiD0oFCOz6sT2xehdgYEN19/gTz1q8XhSrV8cKVb6KciPkJL+hyllA0IOMiKek+jw
30gEkDEgexTwbZi2L5cth0yodUuYio/5vThHGAWYNw8ZnftzKzxRuZ6DE3L1MyUerYNR9hhB7Okl
/mDmNFVLiH1h9fP6mytu7CiAX6pB7Zyp9rZlazjwf73pX0ynbpyD4uIVuhQ0luVHiKNPl87S8bjW
RsHmj/DBvk950QxbOaIBLl7m/FMsWfOonHHas7drC3nF35pawcaY5TQHzjjHpidGBjyXlTs2pY4a
M5gRPO+4MGvN998QDLW6F1W/wVlmVDeLYur5IqDUvXUlWffZ3wZ5dmuHTyDMGFTRenSAvJZu8QcH
0pd4slhv/133dZKDTj9jqlWIfjr1IpAwzakCfrS6eCaUILQ0LIsvqKQCvusaK4nQbAzTMk4b3t/K
qVVkpFaDdNrCqwdbJiF6Zs/QYuuZ9qfYxMKulySmPN7urta9vjNlFhDRLS/N+Qj7FBOlUrxf5G89
QDAfUKH/1l56WKJcvSIahI+R8lIudGeidnlu+SrOI1NIKWUDnC2XAwMmNX7K1OibZ77lX0pnMUcC
exctjxmG+yfE8Pgek7a0gWojWXnTwV7ZcTzRafF+WePpHnHoBCHssjL5L/iNNwpYdNkWUnNUiIDl
fuddEtwCV5IRcoXztNp5f0WQGApFvPwlAPtE9qA3oYtnBxYd8ZS65G3fHIebow4GQCRZF+UC15Nl
w0h8ezkzHPPvpgUyPjxlNSN0A/NvIPh0Wa/eq4UELmNhAyQyZgUW+35w9fPYsc6Z4vtOUniBFjFd
tfYKYn2+a5GCQlpPhFIBsnyBJry/Oj9sPkqif/ywe8X5FcuFYcQU8xiH3zkLzL0jokgHnz5BZNlU
8iQeYJ3f49KNYG/eE5oxwpZghNCMgIGyTYQ+6P4TnEmrUNPDIVsG/jFBElqcW9SZ4tlw7Iz9q+XT
KFhgrikF95ZLA8eqIY3q6pq++MEa2tRHkEwCFoUbCaA+dVX912j/kh2dr3RQGW1Pflp+QsyRsGDE
5L9n9QY2WX66MVkp0TNtdtkkzyeXJKaf7jVWt0/PLZABe9XGZaunIbNnEDLJ6QBbb7vzFur86Nrb
Lmevn3C/GVn5Umh2sgwo4BggGAZOLWyFE9nChuoX2v5ItJyB78cMDT1EJF+j8aXxSuUN2CGCeaJ8
Y8cnmE4Ub3vx8nLTSilS2nFmBUMtV9AvtpKke6JLAwf4U7k8Zqj+DJxGQH4jqSpD7onGdOiMYlYi
un+8BO834tDO4ZVJV+BC8jT4Q8FtdXYr2nXgAHvei9+Fiyt0cTkUlbZqvp/Unrce296D8U//PLT5
QAo1f2aX97APnJoTINoGmF4muyHxltWc5KxVaiCPIITSoD6hT08Gz57NNARwUk+jL3szytHpvNCj
hF6g/m2Lt5VlGXPfCs1VV4JxZ/s6bZVlWPh8rrBhY/FGL9A4UOYfwWiL9A9pUEMb6kTYWASCmkJk
Qkqrd1McTPaRwrRWJa28haQYF0YTLABR9emtmJFxapopWOZZOSBWykGaDtQo3t52DZoJi8DdLV45
qqYPc4zWV+GW2LAWVyiyXlK90Hn2xZQJrv33x2qbUYwxwEQJG1bg206j1a1rTgPOrPog0wZl2Uch
iCyc02jvNy90h59/aHhsD+WdfqjT9Rn4L/oIEtrmPFteknT1BR+KoDu/wNd3G4iMnuUrnmgJcq3O
osPBfSSegmQPaCY9DJMAEulGapTiMEeJEdz69oXqV41SfCrMxByFWK+jR87a7F4BGQg1gFzEdaQ5
awI7S6v7J9C/LpX7Eii1jg2qeYE5S71mLDOxixv78D/qFq6YMegm1+CiHG6SIsJEd1DvFm/fiQck
PAFxLSsENOJZquGgYahAd+pn51eQ3ecJMJAVLnXqYpmdUhdXnht7amMgWzn/dbN2LSFqmPkoanxk
TQE5UUPxW6O8lsMZXEGzlTg8mnk8F2kSqvrG18ME6j2XISnpzos/Kkm5BdNrx/ehns5uqh5OU5B9
bA3IvEhVtiGIP0T19fOl1K/90DzU+U+KH+7WVYK/S5ZhLggYM3VHj6pfB91yn9Xq6XbpSriSmsWj
w0AaLj+Ipe8PbLS5pSG1nh1gaMXRt0Sh+cf2I2nkw1kZ8JkXHQzzGLQcA/Kkn6hI57owl4VkEEfH
xT8kLqa83tWGYSd0CKQ4NQBEEPNSod5XQLZd5yhsKNjTrNzDZmWZHRIbtHTpR2hMbsNFVjPyGvsb
usMMUWU6FgJV5BAUoeIbOdBnKD9MxuzrarUYCByqxhWMgjkBZ5QVKd/7YCaKcN0jLuOzDZRui0KE
T3YMU7gYYsYYMUnD63SDRNWwzc0X+aKUmxBHmwuTi8fXqq6U9MjLbz1Xj/jDhGIwMHUk2zUHP3Ae
8v0yOr/XwfZN4he2Oh9MW1MDIYymK3k/L1K3iuquLg/q3hVU000K/dgUKLbx68fQ1yZqDdgvnb4h
8O6D6HTPFQXj34Vp5ykSbhK7txY0Pz6cOWvgQ+iKe30O7U1haFltz7En6gaiYaZxYtg3n2z3h82E
wUxbgy8JJcS0Bv4JanjnOrTs9zvsgYx4eiaMI3r8j6pYHvjSl0t6v1teeLmnARDdNtANlivE5pO9
M0f5NCezQqx35R4aK9ZH9L03liCnwbCp2FmTTn9JyVIwgWSo8uM2AX4IQSPXXA1jk/4kMaYst/Y+
WBdhCeub2kYWUgd6l2ff5uXQ6/d5nhR44lNzT/SGni2wJzt9O04X+HA24uzK6njDdmDxGEeRJYGo
Atd85RjC2K64Rxc0rFQhKN6HC7561nUQCIbFMi0yZFHXF0/RJgY+7RN+NTKJjkDlQremdoeK5Uhk
nzwwG6aTUkQolfCTRrh9A+4zha/G+y7FlPl2UsmLSZC94Nw58MNd1eacvjSxkF09x/KT4B4rVhqw
EDUTdKoeBsmkuvL5cPFzj+jVrIx4QngTJ9xIHljlbKcrj9eW4wpmpAwlEjoFwtINf2Sn7W7HYKBS
kObmsf498CnztHeCEx4lq9tEk8eu3VLx5bZXkxnUlKO3i1U3g812X8P//iqqPgYm+fABXGPYLZ2+
dk1ofU8CKUom23Ck6Djod3tcIM2x012EAT4blSrDtzjRaOI/2mv6A7+oZxRJRctKNh+/Wxr5MiF7
LrPK0fT/No5/MevJxvugG7an3BFKQmcc6deE23vp+Y2vtbd5nmpwXizxxPxg6Y884i5kKwTxSKnL
ggyExCgwtbO+SrYjdFY/vKJWfEwV/XVeia1881PXrvH5PhkZ38+3M0Z2ayy0aEbbBAzJesgn7KEY
qq/6PRy0pXbhtfWQpPdU+swtc8Yoix6uBw1sIwLhdwEQj+meEgHd8o/9GXtyU0DjK4UULBuPcMfm
3K+Ltz3jt/WAWOBhbXJPtlmaVy3iwGuS1ZHWUse6K0EhJ0n3k4m9S5JhdBRwTUHypuNO053YgBur
ZeELQ+1CX5KUP5zcAmZUQYVlVsDK9fJDgZD+i3eHiTL/H3WuAivE8yg+7TZPpmkkPF4jtel3BS0d
QhUIvXJh6sycfM8UORo5vvLPXFKJ+0NuosTVeKa9YCO9dRST/4Wqb9qRNwPlH655NzyvnGFeS6EY
U5DXgGOHTSHLW2ipar0lZwbXdv2+1vl5PnuJlJrAGHQWN8UdH8lbvZyGFsP7ZOgxPEnj8WYYNMm4
b+ZNxgAibZ0N0apxNlKXNg1QKi5zklfEVmS4xYLFmVPmp/NYa3I1UMc4fMMMCzQ0uw1IhvyTSlf7
9+nqvNSUOXf5BXu0TJZ/bRJaKFXHTli4UXBWqBahqx7sh0+crHrSK3gtWEjond7lkf0IBLwF43S9
zqWS4h0/Km2m5j1AHgf5vFjzuN/Iu3Md1GSNVJQnaP/eMz/KWbSAqat4r/w2g5QwEPYSB77wEUou
2+goFWrKBhTG77yyTAcPuuXc+id/c3eyRzC0VRmipBOpveLdVkF1E2DENZ56beIEqogfe6rRiCpN
srVVbpXuVxz49p/gmZJl4jXtJ+R5Aotbf8yLfQBCzdU8BivU8I2rBskx2f/hp5qxez7PIV8izeqL
vx5sncvR8OQaXEq3M5xByGOQW+7ktMQXf7/XdcUGYxbvLRHHYAG5RjMBJeJ0dGOjMQR5i4AzKYGV
ZgySkaEL6htuRQ/Ejm7YqPPY2ZabSqMcBTfprIIObue7coABoTDdccVBaJolfSPwo3kHaJEIb513
EmVpfRzBS8XfYxfrI06FrQD4Rq2wKaBFZIyTUnj1Hh8jnCpZ20eqVt8w4+2ud/w/sBzFslfdzHi6
qgklgMXkkay2amboYs+r6y0trFpS+8QWt2Xy4MzpLHymWOGQYuTJ9dpi0n+l2gLDIqbgImpBbX/B
QIcNuxW75bIVLP6UUqeiAa+4vYMFmQcgJInoceOVTXJ0ZWLka/CuCsRcrJfKlpPbybCbi0h1DGz7
PRDjpU4a89gnVqD/di85hD2a0Am4b2JSTM2fdFPl9Q4bHXzvYuYZ1mZg6F7Ph1sOYsruQJ4N+Iuh
48q0MDdfsfM/hEIEVK5FW7T1Dkz6Ha4Gv43/qYI2YksuHD9dX1TMfkuSZEDQ+4Yp1wyHhEh+okdQ
Ogeks+R0Fwb186f5PM4C8XVDsqlgt0FtRb5+W6EmVab2y74UGfnYVS0YdFnAB3AMvwJ1HZy0sDZU
EI4v7vkNcnisNxNwxcqVKR3zd0//xtzZ+GH3O0fiFLGq9KhozfAqme1L+jtw5AkWs1BLnjfuE1IG
B0+u7RSGXQId2zfDJhLE+Q7qg5tCc3jI5F3L40V3U3PwpVwYbRdwx09fq8qFnfjRE6yoxVYRG2mG
RwbBx/BSTCbd8eKFnCYf/tll6glf8CQvvTZKuTl2sDy7lemqK6gHIRM0aZApSaOV2jFYIgHq/Fxb
eOKAuvVrIlP+ejaWKVS2tRZpLfCV67aAI9z5A+3ThP9JvtyhHioCqam+gFU13heZUWDf9M4ae8Fo
UA0rqIsP89tmOCt0rCMdYlBPrGmxmYn/cj1MOMe2n1pSbBmukB0htc6YOpPtS/N9j93Jyu51JM5L
gObmpyOGdoyUTS/h2oHayXGh3ijyuVxtWVUBQGzNrbKcwrVshgdPtLQ52pcrLlqk64SE/zGSVG1C
L/EBA3ewEgzchbcS252mi5Bus9DIYmuJqr8x0XzKei7jftyu+B4g6Mlp8gmJX0VNOkvYj47hg5n2
3WPyJ4KK0itFx6CofMpXsN80qjR6ID8O7EHM3hkRC6ScLEI2s9Q70yoM8t1kWwyByGn8q5tIwOyu
xAmLPJJHsf3WlaxGBOj3kXGETaqqAY3sKJhI0eKaneKlUhM52yjjzWx7tPRIHA2ObudnGdeJ7rzJ
L9+sCHDv1Mx9yBANhHLkFmCVlV9vm48Z9mcbwScaDYPRy/bZ5ONi5mrcLTSEggJBVGcYr42l8l9P
ZbwNskI+22PxZQsiLlZ6fi9pE+yGI+yuIEMjdCbUxSBlckSxK/5MVzEFBTwFGffS7O0YqYrZePnq
33VCdne/voqqNaB5uOf8HGwweBfEm61Ar4g7wGfAz6G2roOU+L1YqEB0nWqtvtrB/szZJYB2Qj1D
gOL7xS7EDFztEvKHHoKKAsl0279r4syJ2LfHxR+qFVDGsaMya/Fwa2P6mKxRPHotv4cI+7vy1vo0
cPn2MH6ryOhxU2Mzi3rDYVKjknVaBKo07Kfmj4RzwreM2C6CG7zYM7YJnYjsINCcEWTDEJ2l/74n
Rtgjr/RUXvd7q3mel5gcvDPby1qZfGlB0qOxZVYDOposnxQN9+IGCK5vsNi0IfMa0kHop+eEi1k/
6Pc8TslrVd7954edkMk2hfr6vEnTSaUivcNvEpcoYe5uKC/vW8RLrbHCA69JOvbK8fjn5gk40eYf
dSVvA6qR0826CJnKIMr8Gy62solAxf/flDy2LM2Cc0RqTxFedeS+9/qxEc1P7Yy6HFi86TEa1tca
L2p8po0/tXCDo4gW24RRO242kj9Ll7gdnKHFAkFCsG9XvIsC8NhITh6+qHooTQKzb9pVqeoAuesi
Sid0HTZnJRZujZ05Y/BeSlnpdgjw8pcjg5zBOGg7NVOBdR3qBXzbf/8seAyQ0Y0NYnnyN85joweE
2nrMF/uZFrsEzZ94eK9nTMvEh8WXBjm7z95JFceR9SHoJbHOJqYoBQTAOsbgTl2S0J1cK/6xncmu
12ziAbRMC3YL2n3ZbxWrFOHzBhRUhw1Vb8MAPJwF9O9J7vCNbSE9uC+0rnFciMEl3ay4PALp/2PC
KZhRiayvEnvoiN6SG+J66GNKvAoaX8fnsGinOiaONnvIUJxpHeCXn1f+V/RioCxaQ4b1YRD3ErHK
7G2rCwP+QCJrY01cLDS9gO8b8fORjb+EMsgbP7ZAydYr7ndjkE0F04h48bprHreAt2/XXaosGTpj
uQp+4z3c0h9b9s+LDiTvnw6tWZFoRa08yS0xMOp0xWyp3i5fbeW/Ozn62BI22EE7xioXSnm6ae+7
IVINOHotJ+xMBNS+55eE010TDEVOShYvEN5QrJaPmZpYy1fMEqGvz7fg2NkHTDUxyY+l9dqjp5kC
vkrNoDTSQTukPNCQ9LWcOveY9HZE3iOtKOYPKwNSL5bPTCFaFKMC8Vlv5CYB4jHAV99/lD/jeHxR
FOXUVPahjHGfp/JNjYqcbdCHRgxzj9U+TWkMaRs56adx8uTewF25sCrUT6wYp3tJyXwZDSKfVSp3
mCh2r73IE9umG+f5o8WuASuyUMX6ImVtkQ2AdIz4MwU3D9SEGiON2je+1YqH8ag7e1A65sehZ8e2
dAuGDNRvGz0j92v+lSuRRy19Q3ESpYEBfDh3jNPm1GUAA5dAtRcGXBP04EXDBu+UD+lvjvzc5tF0
b39/Hj0hWVRe+F1cHt11dZyATwGGvGVJBtPe2jsamjmxQt/3ZeHFIR32nHSDNJH5rO2q74fLY5dQ
N3zw8YaEv83yB+d2bG/1KuCbMN8z/hrSIoBBAZXnnbkSSs1jgPJoJ2m9KE3xoOB1NFcW6qcDyAvX
rLQAG9b3BqYq6AM0adgAmeRfibQz2odIZPlzIkHDTAYNIRe2Sw6z0zN3uynpYukOVYGvA+wFQWuT
uXxP/9TJOiJk+HbkJV/e6mAOMI7zudKL6a1laCiAjO4AvA22E5XvoQ2l3nqvMAJxl+wwDh2h02Lb
XZk7tbjAUqSFd2m8CCN/YyVGXavu8+Mb6o9JsGJNnd1TQxO1OvKGY6qWwbIEj+PF1YoACNg5/Aw6
ReZq1dbf1JVkL3krJp3NJOqXQ0xAIw8bWwXPvbBqS2hrGv4gy7+J+eBWpJ2yjijfSaDx2YIe9nuY
zi3wZwKZRZnE+w42uhilVHYANgFpwSb4ZIx3+H0bvqMcQdMfMOiBi61zsoRc3aZ/8Cj0xn5Ea6N1
yK4810NN/aiMCCRqSIGEZVXLb6g15SP8/wLvxqItxY6CeIcD7ttjKNv1hxH51aHLnU5chT2ZCX02
tXV/DR03EMANp3LhW9zhe11v3NSEllCmdPBKV+Bg70SXFGGba1MrG35ORVqwDDqJlq7mTmO1GcuN
Cfs0xUkBEK0M4xQkGNd7rQb+uvps6TjExIjlFVsX4qm5XKh3cJL9tj2t119N30cxiQP+KKT24I1x
3UErct6GU14xRa8vY5R8B+2TnacGdAv48BvU2zebre2MTIbWx67bF6hZFUaUk0P96BKjtpcxn6eL
T4lptJ/3SLlUoq9bOSj78gHpgKpA/KOA3dzsLS+dLOGPSpzOzci0P+VvGpyrMl3sIjqeDSujQcAk
D3JcowYh4WSPx9o+3oCz9ytmHRJcbd5ALHWBhF9dcGJV4AkBODFcah6Oqb+IwtbTX/+v/RHVE+y5
l08jyIphT+oTjcl8w1nqAyfsAr42ASxLOEQvdaUKxdbUYH/xiY2sTjUp5gKXkW4PZCOHotkpZNcs
2ya0Mww6oIlb9/KlPK2G2HjhaOdO7yWrg1LoYudRXCtZ12VqMRrjh/bC9cNMwDHc74fieT3UqEBV
8HEL7YrFEr+zP3Gr6my+6k2r74CJdkSTOk/1vaSgZHI9RWQ2xH2wO5We/oK09jxE3gcPSjtuIoZo
1rLUyAp2vsQlnc+ZBc/zVnSVnPFydz2/z6OVz44XtQCPpVP6H/HjLLIm5RQ3WyTBvHGrFtz2c1dS
b+mw4DbrUQl2ObHgdvJLx6dwVBrHJxLvh2nn1z/x5DDCL5d1ZpXRL2CG+qsmYVLNyLAC0mpnLppV
mREJYWzXnazSVqt7E5a29uf1m/EaC/zySFvgQDBcinJkwmO2w0FuoZ+zYDYy1GYhOwahuaZ6oXdZ
4sGMoWPQ8z734gCRejxVpd9sZGIqmBzw7n6vpeeiZ4zjuvHzGjbGMeSM2YUmknaElTW2GAtO1H+v
PPyllnwu8RpYFEO2G2jT7g6aeCNhqWzrmatMI83klcbeEE5chajdKrpz4EKUCi8pracmhqc5MbrZ
PN9Z+knEy/xu9npTicAQuPuI5lrFiMsGwhMEdOTfUmhF65ySNF9YFO87spgyTijbRXHxiiOjNefw
Xs+IlStWYj2IiesGwoeenDUPXHWddjy8LZovcdOTZWJBtmCVi/mMHVs+4W1yzRZm9guGGlaU8VPt
XnBiBISZZ6qB2ZXOOvHIcTrjSWsR5+bmEwxB3U81H3Ggwk1ExnxD9UIrKy/40dq23HujhdgVdwR2
5JTWD7ETbKWTQFG2H2yPab8a9da5o8SrCLPMkgVhM7KyR1c3d/ZN2Bhe88jH+OQeK/Ru40fGwJBU
yXTe3APnv43qIVsCjcarRKGfP3POe2ZmM3Hl5oJ+itBfm3/qSk7pSkK3lEOBM1kvFEOllzwuzOgB
Cqq6p40cgVi0A54yoMacxDpa+igTLIbm35ch+bsxFsnpbuFjWRbWx6dW1ZmGvYsULkvxN8yfXasM
vDKc8bltl7uniFwwPzJLsgeumLf/2yoBlYkIuJ5R6KnVSxES73VpSgE+OwnsmgflO+IB3Hg9sqlT
jRu+vYer9oENvIMwR6gglLRjNHvHJILEijOTaPpMMwUPRO9KPMonk6vJZ/iosUtWkiiC3GiJp2sq
iPCsqHjFfVJ+M9WgakiFEVZnGHayeFwB0OERguHjSfgGPRefaJPxaCDsxsu0i1eXX75gc1HECTRx
R8mks6TyYZsTy+0inmHCV93J0hZKX1cle+YPO0aN9vSkU12tQ8CghTUbouNIXhky+Hnsu15WmCaY
dJmzbmd8u6WkNcbcpnYZ/Qr+qnRoTCYL9sSas59pqwoHeE6s9K9tSQMr64Ly5ZMYLRky5SIuv2j4
P0GtZXjtUVZTJKUJfhQk4pmXM9ldS8P26yBZ5nekbfimmtJpMRbG52vWPe4t/i2QyiqvPlOM5jk/
YGVmeV2pzUJIhGfQ9qQ3TRY0P9lkhbLvMwCdnrDwO2ENbU+j1qWRV0pI4kYKMv4brqdn2JNwIRDm
CMbDsIrvV3RInq6e9rOqkcLEPlU1Ien+1qDh2wWhzlDljwrYdeQ/i7oaBCiBRRltsKEwkeE6QRD/
zODFO8yEG/IY99iyyyJQ4pp06rWvi++jZe0zuqxd0xHMk1iWKYL7DAb8x9Kg9UR0/CzCShLSOCxy
7fWDzexPb1k6Xgw/y8q7JbKV7QD+YTnGzxuM++SkUvTs7ayB3cadR14+ZbtHdlcIIYuVSnCScc4S
bHJ2cibHKyUBom+cW7m/9I99foZm6afty0nJ+p2PjjLMJC0yFNnpW3zGYKObU+4TGrPcSGCOWCUk
7nGrDLqCRn1SSQ/2tFbkHfLPB8e2uX9srcnMp5kHhInYFmz5GMrBt03HmvuYnPc+yS/RoMmK7QDs
mbR2zcS+K8ec/M6RxKSWWRruiLGRXJ1KoVcNYYpFtAj2v9URdPhpUiiy+jHkvdhaEZTHq/0zPxsJ
fgT7r36DCmwF7i3G5st+GmmemRd5r/sl7rEywWn5QjLVpWTy3bEY2tFtbrV4vGEnmda0AogN0pjo
DHQpViiefM5CyhoeWg5N/j9rCK8HgRoAp0R6fN/bwKG6gYMowONUrCGRZ/ANJGrbplF85NU65vDQ
o7libNxlFrvQvIbD8xsy/futzwoFwLbUlmgiCbmEBiPZ/BAtI/LblAWxX6xRd0oyFDoh+hfzqTLd
bFms+Not1KaDq1f/1s7b/ZFNwR8pVuN6OkEtrPT4srHR8hm46lw6Ad3zaj+LcK50yEzelCFMjsQT
AzIZcnmLceMkpnMmOK6h14qBuKLSp+lx3ZIpzWSm4EVfs7XQlQkU5SFvlgF+TvFCNqP2eRv5pTHQ
ha3UPTFxCzjRkatU8Q01jD5LgHER9sjlCZsleKz7rbVZX/lCyFGd0DdPFWorQZAzrLDAXmeb+mf6
5Wu5WbucMT1MwOxRZ9g6IrbZ9kTaY6OBFOwTChJa5MVyJQIp1VQM4i3m4p2CJIip6Vy8VvDCCkjL
JD2L1o36VmhxLDfmy4MYiwAL5uxN2SgrilaNT6Sj7Bibkh4fBpymB0xitg+df9xsmtgtimIVLOJR
HNfzJ8hQbiO/JhjVlqfjAXQDU48+KbePUuAgF16qpM+5BDPiJ2ToxU9ZjzbYm2TjDMAd7BK0VRx5
aeyqGKrGHKfisZM/cZHAK5C1FcycwkvJrV2qQv8CDcpJpUgaOaz+0vuuyyOVW3vXGZSh9FbGmwTG
EMboSE3SwUUiz1uMqpLkFPh21CjPdkqep9I2aVKoPYNgdHzY+4GgaPmMMM/x67+mDtf+XGUk0Wlh
s3BZ59mUIhyHads477IYgMPkYOlgWsnhJdnt0uN/9/WJTY5W/qSV8TIDFtqIEUGd1rsKwLEpUqBM
6llTODkO5SS0YAbHUNaOJyXZAewjZq/Q4nRB4KzWcEN9LGS13uPH716eKGRzBpe0k8a1X5o2U1e3
NveRAtoPYyowy3eSqiWO+QX48i8SSWPYJ795URTkJp2p2xQCc2yRBoGb9iJRBr6CsqxsrEwJ9Iv/
5pcQwAPQttBnuxuKk/+PRFTKujJwTJdWJOllHWYesJGQDurv1Im8godaXr1ubcxmcb3gTiwCmdH/
VTwFtCqpF2aQoRkm0fedHDObJnhV9aCpTiEoWmVlqvdvj+1Xh4w2Nd6MV2hD+Q2yX4Vsz/FsPGvB
CAFTvXyyx0M1aYixBeLkgMaHscvVX7Jm75VZtLJcy/kJAxt8OEdNSvXJa56rdmvioGJWK82Xjzf2
YcicYUTLSV+fMTjrg+pRpBwiaO6hQ6r4l28PxE6W1nhDvbl1HN2lTxn0zA1FtkCWCn/KAToBGiTK
hi7HuVJ/LPmgIoLCE67iuZE6iVgeXLlExNExAxSYUuTzFtN8c6Zjl9OtvFLiL92m3nFIdcjQ/xs3
FDmB3ZpHv3+OuTTTmELXmIgvDY5afddM27AphKkkMgmwZAqOe51P6cdifqXuYc7d4JVabZ8sE1b7
GFVyjKxh3Wvmg8RrHp7i+Ybo+JZ+Q5qJlSDzbCvx1oIHT2cXdz//vJc4WiW0S+ywOfFHmzOQw/Vi
V55t92LPuiwbBVzuyIiY7DC00ls4WPC+4dDe5yb9NxAZm06FAip3e4eP7L+jBOtEQtGtpvKvqRnO
2CGaULnlHeta7E8E4R+EnaLtRPe1YoKeKXnMChhbMrsS15TJTMvb1nEPVqyQDgaC6l20c9yshxZH
d6D1fZcF8iB/vo3qiYMB/ojCMREcfIpEkT3FkH0qhR2If2DMR5o9SoUfi72pKsEHSB7DJSUmktoo
94Ae2+gyVthZq5UbMJYP+ZiY1/q85+506554PfjnivRryZFUddyis05bCS6E5v/LbsuW0riY7pCz
FWfuKGpHtqJ0QJrrL/n4PW/i4ifSIvLR7/EqJwKbr3eLocX07P8Ai1mSRO6FE5LEfjvvtjeL4MTp
msuXPCP2TIzLDuUnwfB3pJAjcOteeLAXtwZRDbUZm45E1Cw2oMPyqiRPk9p+D5/5wFvjm7XLZ/kK
O/suRK/qHVDIa9bHREg5B3TDL383DuBpY51BJPhv1BfFAXS6nQZSasu2Y2jEr5sY5TjUqqzs2K3j
IWOEVpQUB0KUqEQvxMr3+Blp4rKHyoZ/VPcf1jYvNTHJU1emdOc5h5j3qYynUKXdukUR3DZN10fD
T5ai2CrajXtuHxdymcUSmzWUyDXj48iDRYeeudWKtlq6g+brGuXG1/uL5XKvWoP8j6Ai+2wnoeC3
qFe6nmm4I9mcwsboamcAjODKkafwtE/na70ZTm4+XG+AStk9iTQa38WHUmbyb1JpudmXVGHIurtf
RpAe+NYx13pp2VaMWw+1Q6pl44L/+c9coC4J0TqZsEJitVtlTJMpAuZZUiu7uHadN5blybhBUM1b
mSKgIWsZSJZ4q5I9DQDMPVzyQ7wGVJvZxx53/QPspRKX13rSc0FzM1nLqM1GYpJQ8GLPZf9aCkS6
A1+vCQMIlmC6PPtfvcSD0CThyiuuvUZlmMiXufo3YE8TZMu4DKQ1WgMOzZ1gVO9IsjJY2WUsk+O5
/VrqsmynB0VcbR0J1CanzOlIk3JWjvWKOrqwtOxbTzVNlra7zpf6aXSLI9AX+G3xsPktVqwD/lCb
QD/aqIFI4nuyP5wT51FS8N2ZPTJmQSEQQVYTtLmEduE2gYIDp4S0+hieBWE1NN+RkrgWWZRyVj79
XksBVo1YFP2MCvg8XP+hLlxqQ3l5PrmkNKRnua1LA6VBKemvqxE5f+TXDi5EJwnGId5L0kHWeTzf
prTORWwxdUtF90UmkpaaQq1Og+bHT22cYwHOV5LkSowck0/mPsnSDyFg1i7n+99sKyVEsWru4U2X
xDhoJ5ZixuMwnoX0tz1UelJ4j4b48suQQCSKkWug/j4lEAGxZLTfkQZeLj2sw1wngnhh63EcPrUM
Liq0qnI4i1pJUBAagSVoTifec5Jh6h8ND3PAXnrtiFJh55ne771p8sEU5aJuIMg8sVuAM5C0ATkj
sGpcdSHgV+BUX08s+5t/9gezRI1i8PkAnYoqXYRk2UByxAOsmu+Mb+WZ/eBXnW0Yccq6GW5Je7K8
gRokLDOkiMYj+JGXmSuLTZkWAIzKBmtoja168V4wlcj+V0jyqWMMcJRf+IJfE4t6Y0J/nFqNeG2Y
12TXfHnvpE3MwG4dGmGK42ElHB1pDYy0QxzLafVltyv4LtRL+WI0bJbBD4X8Z1foBMgPaSVL8Vcm
mG33rHgXLhdAttK/n85qS9xEoYjKBD1Fbdn77MwdZF/6gZMRzCwuc7mIP7OSNdQB5c+qOkpIQzfH
HVH8d9GkzhxyHCTJdu5OQKcy/cRkObfwZvId0SRivS1o7cbrWL+AygXhxNzE32pL5cPAc8a0X3Vj
IL6fh/OFjMbHrlGp4YNKSqYhDMW1qqyhZPQGwVguifnN4MT0o6QEMJCg3kxf6JpiXLBGlFwi8buG
7FcIjFyU0RGAXaT/6qElGZoTvhQnzUQavf2rUq9Tt2UL4b7i7W8nZGelj2nD8JGN/UVHbE9hkiXq
BTTMwuxYjnua2vR4Lxh6W2DiZquhAL2qvmp1h5PGdjJ4WRKJxJsZS/fbawsa/59+7pwAZWVjS9aR
n7jf6Ha0LsrSggjJR/CUUemjca8O6GZ6q/OrzH1ULGSw37wKqflNBlS9Xr0QXVqEr+uY7ib5JGYN
g26P9y3qX2mqxFSFf4EKOWlBs2QubfftooY94Z01AJOiEC9b2+LC5COHoGqK/MG7KCer/9ynVxGq
lyxHD22mWpN1wDIlXnx/CSwRFVvWz3XjpXZBd5FljYdpOD2VphB0nrf+apAlTtClcunJ3cdhxSLr
IZT7RBqx3lXhoNtFjTncogosMntc1Qd4SUwgA2N0KEuKF2aJ/rury8KfXaHrOVADIhZlNczRRVKE
RYIgXIRwUQ88+URib8hLHCSG/gmtKzYFff7mPbkHkHwO/AOgSAAX1bpoceD44DtJWtmgJ2WRV7Y8
nPbXSTLPG05TSmSGvxpOaPxiNflMJ7A59GGPFhpo1gtdVcPyyOGFPd0Zmv+FDL1K/ZSb95QZAouO
G/7ynpxifPOZ+LkNGkegkG/wl9VlbArj4/xhkA4Gm3vCqRgd7RV9X0HI5V9H9pYZyMaLOFBKjDr6
ozQgy5YRcJcncYctE+vwLl2oSlFg6gO5SywjhlQFki53cQ8/NJ1iLEsxgsdSSgpRocjURU6aruVA
mT1sRHM5hpFW+tZh3OgO1yVkC+6+bLfis32owi+xvzCZjLn08K55uh2eKPvwWF0yzgAvR12kBAWL
byNxqld13AM22gThLsZg20FTO+Q8PHpxTfu4LqDdJMcnBm2pzZCtE9uZ61npa+Mesa5jOSP7KVQa
tddTmXThwWomJj6uITJu3P88vMJyLLzOvLh0Pp6JZ952AJdaczZNXpHNZddUz6WNU0hhYQLD6exG
rGgLmiNyICSQgXpcL0pZqxWoXviHJRbYLzZ+iL8NSB3bQpZpocjWk1ZiMJIzuTkg69D4HZFAuh/w
j9/FylBsciXZOdhMI3lxHotelWBVZ8P+nYEvwHQhpxrm8h2JA6dv36PFvPRwCBl9LT0RZOisZsdP
UC2neHZJ7Y8LegjTyUw9ac8IWYmRy6DWIFB7c5dspAmJRbWQTmxGsDydAzefpv2wGVQhtA1ARjoh
qK3q28jVLE1ib02TQO7hsgDwbknmm2XGlhy/K8nTY4LMvtdFpAaobG2p7foKfcsuuG7q+nA7t3CF
s+S5gqqEDFdSyJYC3RxAJuSA8Bap7OI4vOIhb8RIbwND2sxeQLid6dmevaa4mEUkHvGyL64Nhu7k
S75JqxTF+oCS99/g8KnytwQyMjjRORR64+NfVAE13+tfOWGdfHuJv2tEB7ZXQNFslKbClIlSFVJC
PgRYMOFhB3c6i7iJRqpqx0VFK2/yEADv5DhdISpWSgM+JxzYJtiz76pZRkwY8j29gc5jR1pdMNjB
osPZJy8Bo/awRuJVKkIJvcFXMUcIbpmq3OAz91pi/RVm3CzRhr13WQgFWAuC3GNmBmkgL8K9VsYu
/9XElqSv8SXd5wdz5ka+Yri+OqPMezuuE2IQ1oDLV4lWeiY/FnogiPrjmfMK3KcBT29qPByJ4NwZ
UikYctiDAbZeKSYCNBLyT4jZWdCiiUgJ+W+Y7J5WcFSrtoKetQihwciQoNj3z+jOEGtoCcFIJxBW
YHN9DTeaR1+6Zey06X1/V7HRLs7s9oyZMny4Eulo1dBYBoLEzZSCOcK3O5cMvrR24W0TWJP8i/lB
C3l5Nh2yAE9sZSktxwijE5ZWVuHl9QlUZ11mlKUvN21RMEfa8sWLe+Sx8cnrwc0rni03bXxWZzeY
MzxeH5UNamW79orCRaim2Oe5f75RPXk1w6vg6rcsusZ7gziv3fEkhb/7yDiQ66H6AEWThxGMQEJZ
L1cbe/hnz6gAbom3b9j1RMJf+PsU7bzk5CDGjOExevl4Q9K2P06R/f1zZC77lvm50+I0J/Kv3G4G
LOnvIvWD95OW0lKv0V4kvCr++zmtAcFALXjo+5Bc5OcyMgHFvC3xOUk/+e5VycD2Vq6jnuFnHHPG
1Qj+C/RB5RjQSvQAVrfnc7oot7Cb7fRCeTcDKkQ5RCPnHuFCS5HMLlLmGwytIYI5qjnt/l5YRvF6
SeFc+hKKybAdTeI6wcSWUpL6DmDZo5YKMvPLuOPLaa4vP38wlbwLLkVo6wT3Up2zIWaGhJgAvjt+
Hai2E41S+tS/w+4lFXBAOL5zmLAzZvonw4Mo5hO9purdpiRzR5wYJPRSFee0UdmtjBZXT6jZVnMM
QSJvIDOXmpMkK2/bQ/fBOWdO0VB/OAiZOhqAGoqiB8aXxMBNMqHTrklhfM/CNOz4PByM6xverUhs
r5RLU7X85TmN0KOoQVSkdEr/KsxyyvvihLciNVcfEjr+GN4sLSUWjHZKM4SnJ6LvAHQMLDtetjPL
xqd3Z2HOFQTp0gaKB4+Xw45nLxyh77ShgtdhrsA7naOvfFHTo+lSGAZUtnGlLDyQ3JWhudieHz8a
DzNP2hoGUYFS7wdgp1wXWQyqexDnA98pwrsnF3V8l5/U7YdQi2TE6Ceca1CnSbRQncxFogh8+hLi
Bg03MgHTPoA8HFstinNj2QAG4QjxZTYUkqq1wbJ0gnTpwuJfFFGQbt99G5Ed3Ogxzo5L9u7ZRNV7
8jW+WOtyiyF25hEG0FQu8Ut0vnQyuHz2aqCVubkPZ65NKKwR0bBldTL/rRXSbWtlnMcd/6DMKI76
5zQGY/pSH1AUcyavC+Y81y/xqpwwfeJYNsKopIRQJ85lV7ZqoJqnY3NFZi5E8IRMdabhuRo/mry0
J3XWHWKnEV6+GAKvTeDJdniLeIFeneWa8qVhpeAae0ZEVRixB8rSTlLvjMB3h0WwhWIbiA74qCFm
vpvfu4nOjqIsA6NT8qfHrIYFlabvqcukqwkZzFfY1PldNudEhffcJW6nmYgMmp3pkKB9aT+HHACJ
oAOb/AwPh3jHKDK7+xqiTbUoWOlk6o0W0vdfgfyao5JYIwAQ+tzEgevEiSOFLzdrlahbeQ1lQyZv
tIjSDIsuMQ0pNY7ZFo4Jh32OZEWoWtne0UgBjvlbUVVoByioe2cB8lfXFdN8BM751aichE+c97Ev
ZnFZszXy3ckKlzi9O5UxQEi5HgUgsNd+hd+IXOVPIsfXCZ8KFG1wYQwEiLmvN9KI1d+AB0Mxq0yb
vxpowtPDDiJbTAqzWtp0qYwKsUWV6eUQ0olWcFC/kWj5gBhulyFxquYIgT/3sEpWjCXspkzotlPD
jBqKjAYSSMlRmkjOLMBghJ57BNhjkM64YjmLbXWtX7x6HQLlgFtR4a+0mWzvCl3zvucjWYw13Dt9
59Gmrm+7Q6j+NZw+bK1A5CsiqdKYFCnEdIZpMakRjz9GoLkE5P/RUbvyvRV3iCG8mB/ruhyd40uV
lCjcvsyb9GfPqjJhhtqdlT0m50v3k2qCdZ7l2KH32n9GF/p2a2wP/uCR9WkEe7lZDnNy+zs9G2SS
SqEsTFvUdg93DEJYsvcMVaa1hdbCcCpunAq5iLb2TdlrcNmFDc5oHRTDRPgoxdTkwtv0blfJ0pj2
3Fi0TiyhFnt0b8wkiL7uuUl/vZQ6UotAUMXc1hv1GF0Mdh3boqQhkypZ0o7KVqQg44wjSdoozcY6
w14t5YFMK8NEMoXl7KZkiPFkJLGEIjBMWldUNA3HhvSZAw8CEzX5MTO0OS6fCvjMBNVXMoivLC5d
rJ2aeX+0xJ9soqbrXXOI/OXBjfnWplMMUECS9w+8XQMA8ICvyrc7WP/hUCLtnWKMu8ZVE/oAgiDW
NEgbarLhr71xyZntHhmngAMzHFaH7DnydjtnT3iZtbnrQJdU5LDTX/6R1wtKQ9dyfiBxYJj/VvxK
7p+SUZgO3OfT04cuuOpxPW/cO1tfVewt271Vp7MNmUebqASwS9Bm9I23iT4DeXjj1lab2ZdPKwAk
ZdJ+kjYFX6C8fg4BKwxbrmwgCk8vuQI5P3JI3uL7pvcwkbK5udUa5gFWLLStyanQK1s3ux+ZRbLq
r691+UnRD/knH+TRyEZ/5u5J/fBdmkJ6qnQTKuD6ws4DjweaNdhd0pUZO7NeWWjz+IuXDxEIYJtG
ioqc0VB/69amZByi9rCBmCRwOCnTkMPMbIZ/s52Ongoid77JBDx3ItifToVxXZKgEGq7E18kIuYy
OUgpV1VUuOAD40rmZLgi6LNk7wsvkM06Wb4v7iHsqSwpvEYXJSu4epmIaFGIZUg8UNhCsC9a1gKR
YhhXoCGrm8y3vANqB45na5ba8CQNfXg+8jK0eEjBJvKCIP8xQhUj4NSM/S70Vjd60QrsmsL3UiJW
3mqR+e5Nk/nCLvEKyr28wfs9ZWeYPvnh9mDAE7FFmTQrQa7f5uaslwxGhCqIXdEEoC5h5QsESCUw
oP4cyE/AP93hFtYczUamYAnH6q0VFAcr//Ad3GUC94p3DuUI+Jn3jazGFtPY1WbmHVE3RuBbIm5T
A76zO7lMgQsL41/fcnr4L/3vYf6A7dFEzH5X69zHdEFsmtEaN0TWBDVvGGJFLgjLsl8f11qyYVZh
NnXBuJwe4KpFWKym4NYw+K+/E2rAiwB28gYWDlTCuWmVmXlPbXz5oSPxjuShF3SU0VJIVASIfIM9
HtyxXtLSWU3+qHbx2zGTX0t/5mKWZwbKyDZGIdImxvdRHB9jLqV6Eu5ZRTbfAZZESE+cM1IpLkIV
0TjZLrSO/Rkni7l7x3jGZCq7uILf0tf4IBre86X20NowpM0rlR4bJH/+Jz7Qx91Kq+j5ZnWP9KOx
I3Uliwm/aZlJg4AlF7jTBRArWltxY1EJkNmaQNWvr2+t6nv0G58q+wVZdU9JtqAhKFgIApAqUIBf
8tnKgLe1hesVY9C0gKf7JCKDNCxOdAVsanGFJHncAV6ePGSp17LJgF/KFZSi1cY3zbGb+CvnHfWk
kW4TjQs5rAMouVDfKyHxHT+E9NxadXbrZ70uyZfBm9nCU4EAC7GFtalHL0gjXDdcHXXYp/kWV1w5
/u8IAwCJiB1QoWbJ2DreEjcc8HnOdgEPPvbDWVIJ6esT6GYdl8mDSRn8OHkLKdHRbH8NQh77OSq4
g7dt3fbSAQGpwNSm001xwWILJxnVVzh8cvwPV5tdQdNs9U8fgsQYL0lwEe4Zv9VfRq+sjVFKOrj8
yRR5WqyrPxVAg/tMlFLsaG+aI113/rTdQjpdmqsMK9+RA/J+tx9SHSDCVWxYvSOkMjI971hluyuo
ogHg0FwXhg9cQ2AIPYs4/2OWYFt4MsrD1xvWGDCCkf24bGaYHY3vtnTcYEt8Y/tUzDLsvEYGYc08
1SnXKF7CAadbkfrIDAvMv0cTxkeuBY+0EXoojR2LjQl6zE3h5rWdIBt2iUXsn1QritSRSQ+mLNnk
6TQXTllaWRdOaqS24CPj7JQQlGj1cCwmpuqfMcrOX6AcRDmkbIpf1DVPlBajx3u/dzRrdm9/Sjtl
6XX6JgnrvtSVt5VTLvuaS1WaoRoUDblrwPJRKK8eXmNrC3h8KwcxSUH89asc+r/v4XxMg4NQ/8vr
Y4Q1f3qgnqQEhB2r+ig6O11F+p3FM2ukezXCeEGxWzz1onNc/q3sC/L1/wRKwQcHlN9I5a+OBpvG
0Vn57qmo37xHnCbVZozojqO4QppXQceRB2tBqs3G2lVCe17koEP/H7CYfwEeCKog77C78j6wXzo3
V/FTWhDYXh8NIZM/0MwOq1IWpVYb5k1NjDQ88OdQSw2To6Wm4Yr4OKmYcVCTVEZOcsVpBfwKRwWq
iikvAktov6mLCs+hc2lWiOHFukmtK0yJMa4Zvl01a8ILsdXfsvqJmWL6MC2aypFRTaeMMDEBcdgC
NtXJxqtRvS1IIzAyPQL8sarFBwCg16IqtzyMMDX3glRX+3s+T0Nf6lAywHP5IVid6Lgu5ey4Ozet
BbP+ksWPn0D86aDFjbwWpb8QPh3EollCqvqyEZxVmLY/Kvedb3M5dUCy42/3Gp7d82dFRP95aaTW
kioLUEjHjpgthXNDOZrO6baDZ7bXCuiHrcdYzD0s5P4aQ8T5mOwAEWNW3uWEAsForhiEQnZzbxCA
goa5QgM3fKIcDCkQW4tPcI4kbDHgeXchodctpStENsoVywTEbU4Tbv7CfRGF96wNq2uZWpc4GfrN
AWCXY43wZtAg1iwmzGtpjnzaqDaa4Xg4Wohui2J1/kEkGWOc+A9XGN39Z0mm7JxTe25uECJAEuEU
rFfxMzToaM2XyKKKlrgd5Cn+AqQ79SAz6YaBsodAaZ3oP3dQcjIzVfbMIpFYvDqZIcOLO1i3Q1oE
HyOIh5jxCB3GQz6dJzFza6KA5ORBAj2D2XY3+KNZ/5t0JSto3VHlp5gR2/AITdbxYJ1F0E4aB5pv
sYDKpZaFrVttO3Oqbl2jEDh9od0+p9NrB0tf1agrrDnxVqTwjtaOAbWxyeefnGAEmHe1ocqmftQh
kRGHsCpsyWsF/ReOAvFaOSOfI/Ce4FitBYWZJNIpF4Fy27dHzGruGFqwjcgC+87pfJ4rT03FRu+z
tSuwGokeNhGjFPZwuEYiGCSWEtyP79RqNv/2zMgaHlr772fyQKQn37Gn6lQGtq0jXfF2MyeDCdeQ
2O4F+4tWkGJ1YsZ+2pJF/WPC9a1I0c4boUFKpoDJ/WaS6ITzZFnvFC1e/ucw3t4qyjFpoSuT90yL
69IYG6c+EcaCEx98dyrZbkIdsBLVwOAF1qpiAPp7qFBBjfZHynoLLRHlPXdbyLu69ycGCzBfSrUk
VzouywdBpeKEW5GDTN+gLbJSCHFdG/H0nGoeb72iUZjrIaNgUhDg9SqG+8Dj5iFMXpMsOP2ArPcl
89bL2mfBH4QnvT+FnHgIdL+sgJl3QgsToBQYmwnMKXqgl9p2wKUpkivjk3+4K8eS1MhEBoQrgTSf
hpQGYUFl0yO7oh0MoFOPEZj2/xQcbChWZKyAbRDHsQlpDqvzTzgEkBVxPym7bFMD19Zjy45vsP/P
a+Memtyl9xNRsLyVTrPXGrMQJo+gEkMl9K6rIZU19ijLnfOQmA4t1Biq2DZg11wCB+TNyLp9oZC1
t13RPy8UkkrmLn3SeiNHxvtEK+/SblySf3fMLl0KBfTyxYepfa/dwE6s3TdvQMTQbVy7sw8Urpc9
H2EdJXoEZmYFGORbccEP5wHTzJLWTMoo1N06VrpbsEmDGyXKlw3Mel4ahlwn26yS5THCl1q3VvgX
JOT+e9SdXVPeIc4fuvLncOoqC+0sNgAfL8slvjznlOuCfQfFh+oPb9OybYdlqI2M9z1sRP7JqrHS
WFLWPe4nDQEISc4A0s27k0p3U9mWMJ8oUtW7myIX1LaaUXAxA/HYrU5k5XeS93PlKMRY9gHyrfCG
m93ecE6uwg9Qz+yqWpk12mI/+ED8sZgUQ6jizFQDeYpTmL92jLaeBOp4S3WFv5S3o3yopPm5Svll
jJHp7ZJs/fCmij12WCVBfP5z3CHi9APxSHmNwnhNi4OjSu+YUCOOVbIrLn6lad9k6t0n6mlQWieh
//+3ecxUFdpoFNCQ6MIjIrwKaAmFghoGYuFEJKqajMcCBvxZs3wK1VahBT8qWLfbrS6U6lj8yYZA
RQR0lvtEFyLLDhJn8ynjqcujr0mKIa+y5sq3nbWqHEEdWdU1Atth+1zpwWWplQMawC2OZX5+iShW
Q/YOZFxnf6RDPXzYuQW2Hyu/wk/ncWgDR89UIHPXHg3KOtiO0aEBgPrsjSPRpBHi3wcbsfu1+IZB
H5U+OhYlWYWvlFeZjlC4H72ZvcGtmUQQVoikVJkynWeZhOPw9lAcF7049ZvsEQurcqxSWRW+AIFk
zdKiYPVVhT5Yj6vV/SWq421Du47Ct8kyqNer2CK50u6lTB2Dr4NMNsaaqLfr+rGFrfKneoUCgwGt
epFaeHOfwPP08z3OO3eek10xGv8cChwDhlNIWPBkMlOz2M7w5BD2YZp0KY8kvqWskwFFICssjEFJ
9MnKKgnVjArACpRr5QeYA48ucpsniKZwiFYCCauaDgmSkjUFspBLVec1MDjZfhN07QyOYKY7s7+V
48QYq4DcfWJCXhdr6PYTcc1GI1WhYNrU+2wjs8pt312qdgtMe0GWdLNWnGcjSxjdMA9tpFECgIS9
5utJxiS5qOH/xVTGx7dsllssPCdFyiuIOhxQ5r1pUVGGlmiebZX9bOuRVvFgVi2IcC0QFoEVYTDZ
6NEvGxPHIY5usBRcHYfcDNaQ5Tfafe2iHTLEMF7yUy9pViBxC2q9+bzmJ6SaLB1Al3eu/mx6Vue6
6XzEpHeMska12FIvsbuS/Ju/l39BGLNMZ6fPWDX32oI/oizxzhh/5xp92d7DHdjTQDy63lL3bO0t
MEOsW9Gzj9SALm4njlqbWVNGfKOmcufHzBSLn7q21Y2CkanhhG/6MgEsG0lU40jiHSoxY2D/sexc
Eq5UlkIy3tN/+i2EgGnUtT5AvBGi+FhyT3jSp4w2oJgPB9iJQ+PIp+g/I8IUlXKm/RcnVcqB8T4V
ssymQbLkNI9UAmQhOpAAX94HBXRmGD2oe+AEeLorkH1+9ekTFv+KT++uVwLvFCde8VfVPEXwh+8U
/yepR0t7Q2SpSvExycGDesFcXsH8we7nAjeLpHhG3fr4sMacTD4l31HVGiwUNhm/EAPThTrPowsv
DObp8hPdJLvghrfPpxbevmP3tszPVUYF0hED89R1YBoc/YE/BJb4AejX4oJ/I+6eM8Um+ElgS3PX
EXbEtixld+9MuWUL4c3xMiFEj/tu2fu2l6d0M+typCRQN+NubteaXASG75znhbXtDEYtH5Zr9vsg
vgUfvueUkYsg1YIAPe6AeFOZXD26KlC9UO/eyEW8IxFKrw/pg+foBoTadxhiX4fidSaBau5/I/1N
Xeyp4gUIAxBUKpjrLDWGTiwBYkN+4KKOVBXlqTQE882GJWWN6pKIrRp0KExNoKIl93xar/pbCUqN
/dA57jHrehIt6PtfFTMAS+5u15xFgREZMuBNwv5GeJs+B4leu680SB5GztmZhhKqUJfasRp5RJGQ
IkuMAKaBHk6f9SdOx7p3+8mn5+yoSV9WfAD5zNJQVsFivgT1OxKKVoih+zLdtzRtHSm7q+mlQOqg
amL6mOWNir7hozWR9ei7Q4LEQXOSnr+jKUNA+t7Z944EYf1A+qQx+GrpMOaK/qJYMCakSczuEudV
J9j5PX94lxlLP60Coo3HG0jdKzaurJhIrThYhpV4bLIIJ/fS2rkv8C2bUeu0zL0HKM6eIlh/j2DL
Hoxb0U8pk1TmwjxPyeWAhS5MHVcCnufl89AjoAskbUAYQpSHvpFBY5jw8D5cZAkEJlHm1Otpdx/X
2C0VPnsBVUBsBmfHgFB3VbDhbzRkYcpFVAKCZLX5HcyGeOrsL+txc8m+YW2iJIyRSKtwD7BGIakm
MC9utyPLquKXYBq1PX//WsRKyvflbFSmCTJur67oHuaR3CVno3N6uxm+8zlfRxLQxp34+LOfDbEW
ShQDntS7jXk91LAsK3PnjVYzdzQe2CSJ6MastQW5xAqyCVLdOTI+N5W8UyfsfTbbmQ28A3ILikjp
vKEchfX2h+1YXmovUuuOFV/6XSeI7wS5e5mUh/Dvxsbj0bdaIpdhUm4/e0Vx5LS4RpufsNeCcZd5
C1aFMHIA3EfBY8CRnzkY1XlZyPAWX3G3shCtUuEDqRZ046w1mkAQrsj+vFyAxc/VZyt00oHY7q1p
+EH0OVwRSCSLKanCU0bt9O3RBZEhUgKo1CJjIY4w/17zKwDPK5y/H0gI+Jssr3TkmthwcspKxDMQ
hamuraBZNHmg/qn9QPF100Mc4z/lFGT/C80IoSn0JJwgoCX0VFJL7CKIYWBUKV8ilMN2TJmNDQeR
TKClhQRMV4BYvZ1trCXOaJY8TjHYfJw3tbNFd3pTJWe2XINYcOYkhvntbadvafMcaB1hSN4mDk3I
KRjA2iOQioQUQRWxFwl7/vyhOyI4ktWPnzNppvn3XzYhmzFDPP+1rQsDrzMZr0NjpFhN+8C9BUAm
xaC+Fo4eGK26WgFe1yB1mecSErI6ChOkLG2cCEgv0PmavkZN9FubHSNAIdXFIG3DMXA0wjhkhIwN
HT/R3z6cicUKYJgjyIipHMwuVzCwNUMniuFbLcRnuHN28EJWNlclVZPVoUs9N7dqYyEQuFMhpQLm
4aXRarnf6uAqLF9cErzSMvRXPwdFdJwxqD0rcUSkqRndstvFQWkwD8EKM55ZIuJ1z4QHGHF6cYyv
+POA8pzchSNsQNcjG6yEaLfejJ5JVh07Juti8Yi+OXmBK5ZqRWPunC8TZD7lomq8/w+9nJApf16I
W6xSXWDhpMCvY6OwmtxCX6Wq2EBqqNtq5zoQQz9P6PEsbm5aHBunSGgQUDrk+3aW6e96v/sWBE6a
3g+E7TJQbsEgeslaFanLvm56XIvNi5eABLKLLpT7C7dz/r/9bH6AHm/oN6/Cd/r3m3ePLYwpADI1
cvp+OE0zs8hWO21U3WdgXL1DjO796+23tY6yOvewd8taV8E6l9fjO5ikje6sFe8O9ibP4H79BeuL
ViGuZLqQ0RuDhB0AA5MF1GyL2jUKm9pr80K6ix2QbQJo6LJE+nbwBiNo6BfKNFOjF0rQAD+zOACa
pP+fgvKZzTsROYrt861Gsdk3CQ9vGqzDAM8BRjEXKE1fcp0l8HTeAKMXOQP5EmjcEykfPFrJFNHl
1HxWd/2+fJvzUQCTNW3cFJRAtsyKewnI36YujPUGfi2PJvyCgBLVyxU+BvFYk9xgJmh5998GeHMy
l/1K0NH9P6SYfIxeibRZAXmXEgrD3Nt3uC8aK/xwxl8hLhsLjuSWeIUBCQ8RZhEURufNu8GHNKjI
IL+JBaF6AmKdYY6XiP1iHoESNd4p9KFQ7xOVudmuL2n1bT+hTUAL49N6w1BWJxvyl0yaJdwMj7pm
C/UV59ydOUSHobpwTbV4gPqhVs0HaOtW8I4rPnG2bH3qQJq7053OjMJSqqeLLSlYXkAW9QCwkeRY
44uS1O8DPXZZF5uA4poekm1bYwqnwgGuBgyza2HyRj6IaeDlsM8GgmTGPm4Nmp7LzyTpwr4bC8EI
Y7Zsse8F1vvV02Dv0HROj2dYujTPC85qnAdIQcLcC8Z+HRC0Mf7xIEYuQzZfyk41kDdrT4/maR00
Dsw4cGonkDLBZMB5Fe0FKF2qKGDMjYId3WEavWqLG1zuiI5GU1IChzS8qH2A4oDMDbzTU8K3LF9d
mmp2GyV3B8zyZ4YObiR5Iu+G0qCwLdGeZTaInhiWa54CSqT+zd/55710pN+n7Jv3eSM0rjDHx12i
eoNJTpOcFNEhs8gbfaNph2Mh1skuv/zE0yIka7C1psVfj/eFRn+hx6LLGZmKIpnycTEk2h+Sr6WA
tubazYTbHmox4bv/2Y9PvcYQYHwSNY7MHezpbdjibOJtdk00gJxgn/YSCjdrgnuTTwRJW4iPmyXX
Jq4WP9YN6vlUlDVFbrPLNCFvvuQjk4OD1oR/ZdTLoDRZiXIXolNQiaxMVn9qCxd9TeLP6ay7JExk
o5Mz/YoOgN4BlNN83d9jUQz+cSaf9zsK64Ip/Ut7IVDB8vvYe7Q/GoY4tjd9bvpYcvfT0MMHYfJz
CTrfsAXPWzAXyhwpV7TZdO5b93mx0B79YgfcxrH72gI1GZ3d/GRDtmzjfmJSLgiVxxhaC7cpOpaw
DkSIwrSiBDTm6KP92gdYwFUQ0RPjjKUdcGvJWC/K4edZoqvSnJ6zEulcxLrEPjC8xps9rL4jgyp3
farRKpQcBO82sv/CzF1xxtZ6PbmQJtwGAWTYCVmw/ajLQpInSOzZ8IGmkBxq7KKB4468zvfwKo+r
frpY/15whSUXZX6FddScmb9zpamrmRRZHUJxcGzu/GDE+TwQpJZDy9xuUMWb83B3FjfwbLwmWi93
0gwj0w7JVDAUVopQRRIyMbxX6xfyeNM/xG2e4sqoy2VQ/J8Z/tbW6CslxDkeaGr4yEupuGdkA/PO
IEqXqgvN64NNV4UFmxomqTUaq92IVwieiQ8+Jj95l/sgzqYVNALkch3asne8ngQJ3JghPbmhj9jb
yXTYWowYrZcqstdPMY8Us686Ux29uLf/gAXkLN9EVb2m3hrS9/plRTbz3jZDXPM0/RxUS2w10xsc
igW9rOxygFXPKRBP1pMJk3F7YHyvK0RsCRhtPveYU3+VekFrkIWzQmnK51DNyPimbzliJhUxhKUG
DqsHTQCr6hHj+vcQlZMqjDSUOJj627aeZa1mPRRQURDwbY3SPDlW+vryiaWoCuAO99OGpbuyr60+
klYzJJipSBBFA5wTJDhwslOrvMMP2seDLZykv+5MRrt2Gl/rEp3MiwXPvwNlRqZ86QhwVzffVpOT
BDGxVfY9vnN5DXKrop8+IH8kbsMtxULIP5IR+qGmCYr0wqu45UFWmpDbHbpDCQifZ/m1vnlpU3lj
m2A8dg5ed0N1zChmvobEnCoLGMSAReKt3UKrkkDODOLT5cxPZdkzzyCLQcjAjuVBvsYlQzFRtMUg
DYuaRmK9i7ukf9pBSEhXBn6Ey7Odir/xuM/LFszSmPcV+/ig5T52rXg9BrzqOulRsj+yx+VS3mnV
K2DeMfhVoAcNDh4phc4W6bdIv0Wv6crYPgYOzEKSq8zUbsgl2birNEBseVr/Z4zqz57MDRjbddpL
WUvhVICntmGtalaDzs7/jAUjYBBAheShNgNyibSCyffnumAR80XNMo5lMYB21RotUKEz1wh0gcRC
qkyV8D4tXhNhfUa2r9Z9w86NK9NtvSwjtTzeg9g/VkzGrQ7NZOIyqpLXErcvqjpt4FPX169zjq3B
0X7l1K/lbrLcfca3k7wvkCmKE/9atHyeYHmQIwd6J1vQTx4Wns/A1vTSH6V9VC+C3fhBfLQSDpFi
Et7+JXCpkRho+ldI3l4XhMG26uIs1FdAyaOuMLsALfZlMpFc9lcan480tsZ8LYf+sFJnLprFJAlc
2wicZt5H4cm+cBnteZ4+7w/nUrFK16Hc6ZuaHNNn66RAjtdkF19zkSU0RSCu6dvGswixh/yTg1Fo
aEu+DofBg0wdo6Rcv/B3LgLf5XzAUyHULsXX6T9haWtpEwucr4fkLlwDpu/3hP+//6MavUJFwJ0b
Xnd6e10UCg7yMlcXEFPy4y7C5t1p4rfIp7v9QpspD9K17F5ocvDBHm7GlW3OebHhm4pN9/Czvqkn
IZDrAba4FQ/UujnZnH7IxHl0epZ3cGxPUwb9Ii3YeHzZRBoREZ0/zLsAdPO7D7MHJ5X1eADeGS3G
nGZFznF2cxnVP0IKAr1ubjLELOtTDyAkiF/Zt86xcAQ9ERkxrlXeL98XvCOIt9yu8jd+XZQl+rkp
96hVyTgSJVfl3clReA8Y1PeAMjvn/4rH+dWdsxOU6o6HwlqdfTFhlBfy86dNWnEXnE6LV29C3lWO
pPU+S8nngIZXqkdzwLfzRNZc628DjOOaXOfEgWSKXYe/T0xm7n4dtHD4jOENOitx0UQgjCGFlFKa
aEsDO5ml0BiDY5NUV/sWj47L0bmvwMwEYhH6RtSZwsuApUwJa3nnXnxPciG8Hey4uFzL7Q6sALmW
gGQ3c5yl6g88sueiTIIwXQ+ksJIKSPCdsf3hv4uf7Ek8RHuHNuk5jc6oUNEZv/XqbHBqLRHxHGxO
3dKQtT7x9Zv3TKpggZI+Qsv0wkpEBiA/V2aLIuW1rQYNau/6P5yLVVN4AZ0iQIqBtkmKqm2PW7XN
V8s7BEwyv1vP6nc/LPXYQcpDf/dC5AxDoe+3wsChxMUIxstzz7Bbr80vsMGE7+ax+c+a35RObRHB
2N+LKxA6c6IT3mQvlLPiAO8S3zADssnpO82N8z/jdjw/OXrFZVj6mBIylhYJiEmycd7w2x4M+FHW
lCEoS/z/UFMVCm3S62Ec4X4GauA8j/qCAMZ232O9T4lH5tVSnswXnG7VzynXit+hDeyx4Z9YGZ3h
RBpLQGDTih7yfNGHoNTebOkacMcZsNVNKb7JZWyVRLsL7nFOkXLxFFig6b3znCQs9DOy6F9BjnZ/
Wv+uQ8urM0xMivjDUyZqpllN9kaIHlRmZi4BnjG8dHfmW8fY39czRcsP4mw941NZYPoVTXhAdgPm
R53yBG8OmICBVsN6uJt09TZk45YmEVwdB4AKNUrZfmj0DaWMwMFg0X6RIoDYkWx+XV+p/KBDwuQk
pVgGXJcw14H/TNlRZ2IKSlkX03YwqQrsmmY8akQos6E3PpzqJVX8fYYY7vssItriw005BIPWm4M6
jpDxq1IFWuqG6I30I9fz671zsrlyPlwrfvI6gyIP5IdJ0wb8+ytWnOjBmx1FY8B6SqFNTX389pOf
SXkb/G3y4GM/Hj5U+VBetbSfTyq6wc1wBunyb+/V+CIaLZanbz1KwTf36FVhAdAGSgwpjOOqAHSc
cVIrLrcRapfoEKLnhE9f2eUOkIatpZiy2t0st9uaxKHL9FrJlFW1wazwzvVZvNCu74zAaWUhPMqS
DxmUk2LDpx5kTSSed+bSgqkCP3S8Ryztnb1ZNEJ5HWLNHIEZuRHTwDy0tjfUZVRTtBEaZgNVUVNX
UHXYYYC03YQGRsLFAsQQ7omIOHnAh1z32F7QZfqDGu1sr1+4NVGhgizP0U8Tq7J2uO29Gakpy5ib
YS8D/oVv6wq6/z5DZTHR/MrdNwQ3TSAyuKcn2bamLcmfTCpp6OfwxtcrBVjh2tB1ELXrVoekqFSK
Zsj28AdXiBA4sqsx/0aZXWAjOEoQwHg5SbU7P474HrnP6iTCcfZgEoh9j5tz0FdRZ3/Fv1V3h6Z5
ks4MK7yY7bAllk3S04+Zw3kgGhEB9ZXFQ+dHtUSs6lZOmhs7glTe4k3fy5nRZecpd92Pl5j8XjLV
giZ+YjmvOK8c8oVXzUspbaU9k0bVlekDKPi9uYc/JurPhwxgBAqrqUn+m/M4R0O/voFWupQsNvVd
QFY51/jxj8phk48g2g5CFmbepurfp/uZnTVZkgppCZEt/xdaF5y9zZKm76x1dbkMc4CsnsOAZdRY
OE2KMpdm8U0/h1YXUecJDDHubZFhuulSi9VKfsaGsnxj89Y48kstjALVVPh7wuC72NkBe5q3XGw3
ir/lCK1Qeo2QvDHOuSHHHdhbMV+S0F0FOZ9fiT85OrDXtRSrdwWMLmPD3uGaoHD/+JSJJsg7AKN9
eQBAULGkZB/ohn+1J+WMe5C+OpaUpFwd6wAbfR0l0q/1BXt79IpE7eUl/QSaRVwfRPw2ohlIjoet
hinUWSFKIoC5RerbPSSt/k2ajC9Sb2xmmlS3F/qIDXsktl2kfSFOklrZQM8YhWLXQ1sI/2VXN/zc
0gNfAUx8WCX97KljFErsbaoDvvadCjPAKjV+Dy8z/mrc71T/hJG8u52uYTjFSTdBsAI15cdEp2Lr
l0x1I6x2iT0C1IVgBVhknbKlvNbK0nGCzMa9WXSC+IqxONTwncNgCrRpbzElX2L2BjH3D5r7I4Tw
ypjhgMJ/PO+/gYsvKhnPDeCj4BrildHmN6aMAWaUN7fAORFBu0NtoQt2Gh9263k//rBeILRxzfaV
ZpoDEmddsAx3/t1rr8RryX5gxbFDdlH/qehI3ow+hNCF9ALCiZ1mpJufAGGBrKsM0ceETvjWVkh8
IqAVaiuuqLtkKPIQCwptfxgnnkl0lXByqbsbRUmL131QKLwzJdcvAhkscJyhGHWtehoF9nmfoLYf
fCK1twCzDhKq/V/WaZNVwm2W/vyRVozn3Qqk/U+pifaRiyiYDAOv0QavwVHklECkN4Ob5kwgwNMP
Ux4mkT2PgQml/6xpi8zHL+ST45NgUdDfwYG5QQTGqOUYhForjc8gZqYMPFjemFpg8wNY2JBPvD0i
Jt+Pi5hiGL7XVZSPK0FzUk074U0KKgzwTFdbmDbvhrVeINHi6UHXVKTVH5CuMq4RDDqMXhpJ4VxU
bkKYeEzILUW17tP/t/PzrHtTe1bFNM19XYh4nxwefz64x6yrR5jxkjKufGqvmYK3HY3kEqkaeF7p
ModXezqDVYEs98WR3WdVpgZb85Tt4p0Ka+oDv6a/ur7/46BkW9eOKsngGGafqOR3AoP/XTyjCNt3
NNJRQXnYH5kPhO/MD3xFk2hYZlE3bDNXDp1YqzD+tUwAOn3EOTtzmSgZ7zetY4Mv90bGZn7t+gB/
pkBNhW9kgKr8b97veGUJgYBz2emeRqIjt+4iU/Prm/GduOmzfB+mmL8IaS2la63XTJR69aS7IUVF
eb5snHlPZpKcDtPSbEQsRG1bB8w0SDibOCXHaT5t3Ad+Eb2/af4L60m9WHtvwzts3Ft/i5SUUa37
3w+WoY1haX6hw0HrL/ZQKfIs2QW+tps1a0vQCL2ysmIyQDglHi/i/DK4T/wePg4832MqQ9pdCUDv
dCM2lKWU7MlQFK0CfoQXO1jvmyN6RHnzZURPW+NpRuL2a/o9HWsgVoY7cIsHph96JvoUqO8ZZwxT
x89R+0Eq0AkeoB1nh6o5LZVFi9BV9xuIry7aP30LNUHm06ntqQDZe7X+c1crHskWzwDUAiqttRg5
g/DM9QRFlniJxjMtPub74dwwc1IwMswNfTqCgNZE3ANkDvdfgb0KLwvSm1zLaZyECCkvIswIXBrp
87HCHCPFjgMCTmS16GT2jzseooRT4Ycz0kJ2h/X4suUkO5ZSt6JHh6g5sYy8AeGCbEhK/exAMx2S
1aarsBia9Rw7iGH94tI5D5lQg5FSnRfVfl0nPSDU7ypuI+JRlReZzZQ1ZXW5IEzvn4oxun+2PpO/
dTzXFRhYs+aWPepIadGlQAwrAZhbwYo2nfFYQkzgFMNbRri4wHa1M5wPFwrEt7aEznMcjGJ51kW4
W0AGG4STAkuCtly9yDu03JdYjSd/0DB7BpzxWvFL6DwJmQ06T5vdv22v1V6X3o5566YMFLYEETeH
ORA0B4O4r5BTmnb05oTJqi7QDl+yFVEOX6sbgKi9G9kErHrlx2gzdaI4kD+WdMncJSSerD5OphxI
Swidm/8FEmU0kMsOE0sx24jG/gCTbhtU8VKxMpqyf9/6Pg4XXjcPU1a21i68G20XVnhNgR4ykEER
oECNnpFV3WOkRo5gl3MR+HmoXTLJBLjvtCiaCpOgp9hjKz5MIHWrjsordEFc0yOkTtnDFbNbB7EQ
izH6NWRnuVkYfR8r1RXY93fyzXqrf2cEh2X/whtXn16fWzuPpC+gh82qxh1mo7YmmkiOEEsYw2eZ
jUQFPlrr1nPdv/0nHNrGtFDZVQOG26GbB1Db2rP/RnclFa8oROdB9u3aOHmQrbdsLN+pwdkshfe0
oBlGaI6LP74jMvrO+bdGLtyMRAFBw9DXxsUF6Jh5zKFtMVYEl3C0WacQS0pQW/RX00M6k4Nd+CZk
PZGRAaQsI8F+QagojJyjXxN8gHxorUkBuCrhU6JOprve74OTjAgSt+RpMrsE6eu+R2MFw5f1YBX4
C2BIL2giVYtK/2xbtK0EenlV8Qkn+J8YMwbq6D4LLwabzaqwxudjIRs5pgZoymv+0yqmjaLhD23l
ccRMsgvup48PAQRPlKRFJA10D7E9m0sAo58hQ1BwhWgt22y3hZUl+79wI0r/tIA2BfVLWletavZr
I6YiTtp8PMczj3ZjC1COesuuWGrDE7la5pT5koaIV7RfkGlcbXXxbezspX7hBVxVTqFNAPAna1ay
Qur0h+G0nHSIOiEBLvaYvHJXoOC8/P54f5G3neTrtEELTuX4kRDa6N9HTpnX+We1YEDfy+snfZvy
B1B9+tOjUgUpux1b3uhIFGt97lQIQCSqoMF3QMjHdviSjhHXxQxbDOqNOgfsKU24c809VehgEU8K
0WH5TJnjCtF4vN3dr3WsjEovaMz1qTyvvjjfhzsVHy4gBt6Hd0yCxaiVYUXcdQhOfVdCBWEGoxWJ
6/U3hijTPK+Nk3HPtlgicJtdCWEqCobU+3PX76yHz4acuxv6+lvvnTjslV14nehL9yZNFJu8kJTG
e5ZXMPrXNWMOQYjAVsqH8t+t0biXnfj8qD8/Vy4oSgcp4e1WPf9Ez2SA6XXw4HViIj/wA4J7Fkqe
Bjd0Rd+/XnJ8ZtorbhWCcmagmOkD5wHAXE8xmjtWWuHqDM0+JmhyXArMISfcxzzR0RWQRhn4OgE9
mq7qoDw+gdU29cxEQ1MYIV1WE6HbUE0MX14H0skdJtT9i+BGn0uVM9HAy+8CtG7933wiS9KXMake
Q1COHw2Ipklrbe24AYAdZyiMSfDh/rVDQjcRQHl8X3dIhla3tNYcxz5Djr8HmirY7xW9/hjxgHrE
C1jg9IBFEIUotJOjOW9WxUvsHW9YiSSZaNX9ktrdUU5g+R+QQZYkYdh5AN3o/xC2EVZfSKUIvMjZ
27GHFfVchsrNhHfCaDrevnBSzVkvoV7aBA/G98arTVv8N+xPw733FgnrV47kn6j/KK/XQ7uq63+H
0UDKxuWU7W5VABlPgogzf/IpE6nBFKO7fsDDkaKvQI7DJayCFcEYZr25X76xjD81YcUGiT6vruN/
50Cr98X20ZlpGMejG1rREgcnVJik+3dXVnG+GiZzYaMZRQKLZYSHaRKu3qUwVhg6zf0U7MWW+oHc
bKwWPbclMxYfLoHRPFBjvVTCaxDXfWSqol2rDGWC0f8AiKShXHqqf7YUi+V32A8eqsBzs3Jt3Ju5
bvNM4M2+N0qBwtIcRHistTaR30OgrO1IXzRKax461JB3BmwPglNQCdUrTFYla0uuFVoPWV03F5vU
0LSIfpmOvJZ1q3MUbb/jcGC1vaY0yNRHfJuwAugDKVdU0IwzH5NZ+n3x0mAYavVlfSfxmhvDpUrO
jSFhCYm5EwQrYlqkMWapazPCpjP8KPI4Cn+jjjkx6m+sSJ5EFfX/GjKV/P4TWs6ZjXtvuVzsJVcr
8Qv+dda1xe/qHeW02KmjwpF7s2QHWzzaB2K+lRyYuOKUhrPTAyoJ+uGMtE6g8+N6h9GZn4N/Jd92
Nlut+67UnoRrSJHF7iqP4k76HumyikOmGGH6G8AKe65nC1RXDRj+Fqctd3j02oENTxqba6LvOgBS
VGS3zlRBFbD2MtiEsXscQo/MrSO02TavkTxqHiBiqtk6eTiXfdDDZ5mVhoiBavNuMr6ybDQ/thj1
F99AfZfYLpT73U+HS3y+9vz9fsSXYcF+9jm+XtlC+ATQxHXj7UpYdch9zzNk7i4Hkn3eJgeg40Yl
u6wBiLzsG14VLLVIoGcxP38tzLQo8T6Y81/glhn1qNbVlBKYdUYJPDioUuVyWJ0vt9/V1dK/YODe
i8B6yezRaEUFWAJaHMznJkEMY09GPRI4rgo7shph+1NCAhQYZw/iA3JUZHXiFZZmuzGiF5xWb8Dy
IoLhnpGAeuJL6VjsYRHTh7uXb9yeEyRPZjYCeD/Swie1q4R2rHq5a+9IVNtomUJTQo2LQN+bqRRb
JY3V0tHFqfovIdQrQSalx6kZwj3LkUhvlTSS0CkS9tq1GpI7xhofWPpxcN4VJEw4h649c4ATfZMW
j1qyqqg16rKZRYhooJ9b8Sk4FvoB3OvqliWQBt2lczzHLReJCDVn6DJLGDPZIJoLKx3QbIP5qMiL
+fWOUOLCiKZvzuhZx7Bet9eU0sFQasw5XGIdvojTIi45c3AxLS3aESzyZlQpd3fJzoo1nXXXUXc9
2ApEWUJytN+Z6tc11nvnArN433md7WZjLn+JrNGF/RfX5umaLwObl1GT17PvAkUTpqMtX5ZSruLg
pPZkazl6Q2j7vIOavdHjSWeY97gWiD3jwVL08PJR9iV1VhfD9amRXGf0Z4Lkcp0mkkHgLsvHV4PG
Wa61oSbJnSpKxaqWST5u2sgoG2sGU8cPYEAiwVRY7J83dCSY+em28EJwht25smZv+J49QR+edJyJ
md4aM5OOLwBVmyqLWusT6EDrU+jwfub0evoIHRXoMSZwCRgspS8U+lQ3/XxHpzqx0LJU4Ue8f3MA
DD2JLnz0M7BM+QDOmIAxf6PviIjOhM+R9/go1+Wg4jEfq2/zK1Df+h0Bso7txDxTN7jXaDcujpfP
ZOlTEFEjdedMW3w6Nc5pBKOTn/9bl/NUHlLWBTmImHpaDskrL95uNSsC4Xia9QGkSqQ7blBOLdVm
5+HMbdlDeZ2B9G2xPysAAHjia+J5KzAFq6kvMFGR3G2fbhWSMicfAq+gyIL9dHAO3loYZv3p9XUm
jExgpAef4pUcjjaoEgkq4MiOUEs8YTMy9f8UOCe1X5DUC1eNuaKUpACCTVrINUB2SXRPb08Stlua
1xRO9uSdRZCOxeDsl017kAXlFG6I6OFAZxyXbb2AE3IeU3bHJ4H/eBPZ/VZr/S+DDZfBwgpafAos
HtR8kypVtBQmHBHwDofTQEDVreInCEUoCjqSx+0cUbxXHU3Hca8cVdL3W3pvmgqZ8iMQ2yAYmVt2
SoLHZvWYJD77vQ0RRwqU+QCIO2J2vcTVgQ//Co/0d0HHcpNhayYwB3C7FPbaXDBHr8Dds0ZZlADJ
AurhZCdHIbfZnhbi4Z9+rCh5kK/th0I+JHYXZM2VHDAHcNfHBKKepMomTyhn9+T6k69rvwBBR3A0
oXYz4PBb0oKUv1JEqjMSDsXOB8d90g6Z6kOfmenWc0sYXXzF92y03BK6/6hQ5XQWVPJVE2CnbvS9
l4Nr2C4BvUhbo4iL2HJEEH5HzUC+jgri4O/pWHtTjmMWcKmflnnsxQN6b8Vvts2LrsxY/hCcWJgA
jsLYXuPzirogui6e4S/FjxrmCagUB5WK09P6XpmJBe+Lmqbj7He/eInIud4IVD8rffoXCsMvKqT9
70ZRrsbPRJ5xJedGZyHYzZtjcuKBoweDJgg28v5m/t5utplYMcNZ2WDSP2dRvCSRqr+Um/w3GWqY
z+2u1+NS3xdovg2VMbl1sb8RDtyXWWl37R0RazoKYfwxlIMCNi8j6k49uhFsEcIe9zfhkBMz3vNM
oI9DDD4PGo/XNRb2DaT2SPc+HyvosV3SqlgT9AIJ4+XarQNFWEhoP18zKc+bjYq9oNRoCQsGmlYP
PcEo+UYMSEX6f1culQ3gArpcl7/o8vC13lipfu3IvAqYKPAFGJK2tVFwjE2mLOLHsG7Hd2g0SN+V
OxoY+ZVvDfBnbxGMfblxP+WQkjNIXccCgfWmfM8baI7b9uKycsWWeITWlbVSkLcomH3qJNiR19HG
hmsDoanklfmURsXld2sFxTO8kiqV2Bot+k5T+ozpYgK8oU/Gd0a7gvKoShPGRb57OXPG0sBKVB/2
EA96Bbhcl9U55Rpa/JESo0U9QWLcqvmKy4GeKEQUsWjugmGcoiv3wNYtfbyBGlMcBnU2xKmovk7S
raz7xyP+UqTPEPPnY//zn8r4ENUyahv0aUAPS2ZsB3TNyOzbhnL6ytjpa04dCyuBEL6XEku3tNiB
pSkSzft2G0c3FjjRFw9dIhHiKkN5Z/9KPEX/4TatHTTxTo5qpP/lALBkc1OUxwjuZfVXOEOV53Uq
p4z7ZN8r6Rr3Y+ozgf5xb5RRuSPhZgVYEDu2a3dDdvEsDgQnc7F4nU2hQbpNNDyKy0VibEAKiwJU
OhRAJZn3wmwzD5tv6cQPPnT0IdgiaRFw1rRN7pbXbuBL6JR30OOn7ycxvoCUfUoO/vlREOYgq16N
eUkxghn94OIBstUzTQPCsvi/vLrjXUvZKlQA2iDFhBZADftJLQKtvq6xf1X7HEfo3V8IcWSYf4ht
RyC7lYhHJfedVjVmETwM+8m4B1nvg4XgDVYIWFJilm9eZSu2WispI2Cg4So9h7SW5nWLPx0rvEsW
OfcPMLTBIy1Pagvy/6nCgpFaWQro8ykaxCokdToa3LGe3+nfuo8FOcsfXpRqS9GaWiBcQ1aPOcIy
5bOdVIMlHaZNkC91T0C0OvbY3IpAYp9Y0vcEJ6hjL5PUPJL+eByGWzVXdQ9FGfqwsO9MSH77+9LP
H4fSUi+3LLH0upECcT3l8azLrFt8F6IoucmnQaKq3/vG/7lS7ngKsDvXcXdXTBO2AXPq6y4xw+MG
wlAUUajDwdaQWwGitGk7kwA6hPRnx6TDA95keW2voEm44JLYtXd/yfKXFM031I9TKl8cB46/O6kw
EOkGvEULtVdT10prprdGrlxaXPDP6fnTL0A92rpnciF/mX/3GrMJKrttbfssjH0aBusFhfPWlggn
KiLpFzSpdjclPgdNFG4gAeyTC5MvSjNKV5XNws6f3iFxvr8L919Ufe1qU0igTon1Ol+kEmKkoP7H
rXF1+Ti+p1Vdjp+ncOrBT8FSkJSNdqduiKqAM4gE3ZXQ2tH4395DSyXjTte4WvopDKAMLKutAaVM
362io63526PR/EcIkJvBZ4lSLChRRCKPGgQMRzd7+ds0cKEsoHaT2KW+InADkY1lzYKjnjwdYQoI
fcDdVwNRQc5rI76Dc0qtu8kgc8NidNpK8sFEZhai3sJFWbWCVPD2VmzOSe4rbNC8BrvPBeH/Lqb7
3Fs/fVsxNK3RSg0iAbh7qpLEUrm/45Ggu+y0MlfdMcxKvK9STyKtTN7y0DQOw4KjDY8d3PIYIVxX
2Xglhs18xQczla4gvircVLk/nf/FxkUsLnxpcexBtWqrzvl5VAelaPpNs3HHS/UfN52u8KXgTaYd
1xP3npPdjTPIzXJutliuZiM3R9kq9x+LYB3qJBXUvTuJkEtt1ywbeU20KoomImYnotkKTtA3wAij
JO840nyHIwC7mp39BE5uDpn2RSRsOnV8Tzpj6JaJi9va6R/+Lkz9rl0dmvo5IFLGl4Y86rSi/A5e
qySmokQ5pZrWoSDpWJuI5e9mDAb2Av67i5K011z4BRyeVhTgtpPVodbrEFfgieai8mQedv5eVKdR
5GZ9BMQJvw6gJQmo9yb2XvbQZCGhiVtYj37tIkJEiyNiyAIyaGfvPKFQ1HYZKvFJw94Nq0lAH0xr
nxu/lpV5VJw2t/CA43fVEa0zVKwBNWzCy8t6tAhTU2zjNXoN1nQgOcOF40FKqcmgKvGOW1WyyzLM
E3olO/YNeXAIRNe2BaKfWheMm8e6sLG3gbwMv9QW8F3R06a4+LfNXYmch8rTBc86ou8Jzepw9XNq
8d9NFJXP6+aI+UUGqAtwviqCAWWA/WQawDpE8KfYSMd6eZ/tTOjq7PsCoGAx/2lIuCmkGdNbfATg
+SYa0lrwwfoHNUnZW3bIQ1NcjgOIy7c5zuf35fgkSGNiCXoq263yCX4BDOwP8q3UCBLtvNLAsAex
JxwSbF2Z5gbshKCBipJ7hwTFQOZBX1tDrhqHGogzJy+TngRqf1KmZmcCTKXsG3aFi2RjmbLFVSZU
J1mIXAwsX+1ZxHb17aUtJ3PYWdiPbJjcIGUCgi1jRWcgkm5xTK4wLTTosGTmG4yImA0P7RZdecMB
SQCm3qEItx/W7FU5hftX1Q5+LR3nNVmbghpkFewDOrjRznLohr4WnRqx5CCyeU9Ii8d6zlpLihpv
AmovNjYUUa449qXvDCWhl2BVea1pL3PrnnjuWDQR+FQlCooT4dgB4lR1rHGzpaxtEU30PhPrEupO
ZQhWwN6Og0G92rXUf66GDJju6OI5W8xYK7XhqfgKE7/1ysKUtlfnfPOfb1otZmT+hzyY4C1fvS4l
PA1p0ZvOVGyko9Jf4AZARh6U90WTJmqD5jQQXvOBKkTnqlJ8PV7tffzjpZwT+O0R5iB+K3IxwcrP
Z2iTAYRA0rzjQ17cTBTi+QXzwatgq1rbcfeAR65u6OoF3JnB6SvMb/rD4SLSg1d52E5+y3mDjLQb
9di9+o8zZYV+wcT9mXoO+22KHq05mV5bcHHBsB64GwnBj/lamTyICPqhwpNlhZl8fUfyuhrdeTMO
Dt8o4ynpo04xRlgR64blDABBYIOVPO/pRMo7JEXqDSh8kokFmxcghQmJkw3lME6KkKyyi1GqdE4q
66OQeN+xT+mxZITTpa+CDmw9Gqut+ta2l+YHvc0hxafH3pnEz1PnNG4ZUVHx2TFOwvqoKriVN/tX
fJE9hAOPtn22wHNE27Fa7mn4XK6F6x0+gnr19FrO753LEE86PNQhdzSuSQZpFxvGWgFDShpUxoOH
wDqSBWOtJQ4/HPfErCVxkd1rksw6AbNIUWK77rdpbDGUrgMdIcEW9eA/M91KBOP3rtNSAZ6S9Kpo
SqseOZYn9z4CK9gD6fDXGU7RHiJ07sD+giVGJzV4u5O/GBoKwmus7tqP3+WTf0mNAe1wIG32DjS7
uavEb13i7nGWaAlbhUzQt01o7FNfbYnnSbvKCZ70zgPJbybLnYmcAJQM4HzEnUYcASRc7iqZ+iBz
BGmLw0zCwfy/W309zNYC6n8JD/VOnxCMUg0WvO61msvu3jBv7rUWkehyvJzOFQGNY780aJfCfcpZ
s61GJVoHHIPxLZw7Jdzlzp4/WioUVJ2wy7dVQpWHhdFdkNrXzi7y450iED0ejkeQlUpAIHE38i5T
CRGS/dzRitbD8OVUi+KC1C+Kz7fPKgb2XR9Vla1O9lbrulLwVUQqsqiGr3zp076Oof78u+N80Ohp
aKZ4L7K7Yj1vaWT2dATtVqCGQsZyzGZ/9jJaqTvqtk92rqsn+uAg46hlqQLh1lbjT+s5qLKzFso+
P+X7DI0sm2t29HJ/AZLMJX4RvcgiW9fyxIidG368+2TF0YXmAqFp0S02fn9sfWfVF4e8sfgwUh3+
o0X9KRLeMpgMCFMu7jrUUUewp2hfkxSJHFo6bxOPKS5Fc4m/dSTu/qAjapuj8q1jJl+LqC+vqayY
Iu+NumD4lfIrmMpVVGrbnf2GKWySaYgCMLz5RdjS859AMq9zLBgxXO9kROfglVHXvm8aw0AJZxg0
uEwAkGSMDxWKlXLer5SoyszQk2onR4BtRyJ72UOVBsGK9leuIzvjaDY/jlAFroHVbazdZOnvXmrs
Rr+f9dmZgyShOaGTRRYJfocD0pcU2Z4SaS8eaytQ6E4zDT753466cdt9D34vawVf/g8Qopjw9dEU
Sw2zSEV2lo5XRQhnEKoxzBK3A4qF/LPz5L0Nu3Xt3N1+2KPI7K71ZwqlalvnjbLzR7f3ffSQpHEP
bOO68WUOpDTasjlYg9U1l0bvwpN3BOYaGl6yUYJH8Ji0arStrjNtI3OKr9UYKQP2TbRnHSdM5N+l
fhwoJ7IOhjbzyEQRVw8h18oqtUlZBVUE7IHJU/CHwW9e1prCBYhYkKTyx4awGg9Wsxlio/nTgKIR
qN+NR5GbLqT6HunX2WiTo+altduz2hPQxWX6xXxKcFmp+wflLJs9XMk3/dbQr6rD8464uiy1Q6Dc
S3tdRBSHtC2ePeBqVnQ9agrVV6S9xLH5GRegGCDRQOfxbwXyfQTH+LH8BdiCk8i2qVF0p8DS+QLN
nxJmMqV+Paf2scj5y2hoXWYeoPX1svrAEd4HKM4JNb4Ticaa0Lk4s5BvdcZwZbEbhB2dWJaoiUYS
BHOZYlgwoesdXUEBuCrg9YVO6y+LWapW/mQ+2PvNCihX0RrWl/PRyVXN8oHJgc5L3bc7PtUH/bvP
jWP3rk62gQqhvasIhH/1u0WV7dU9XxeNwmhLccXaU+xSnFbSeP5Tt6rEt3WNB9ey3uzYV8SUOQNL
8rZfpf/B8zb/fRcpnBswoM8s8VJ3z5WvykCs3BBU7avLcyANh1NePnaN6bC1/579ZnKjtw3RTIxQ
ESsy04Jm5zBycoprK+8HMQA9sgxSh6F+IebsJBlNPUFsa6Xl5yDDtYwytyf8s+O4Z1Yntp3GdBZj
3k7Mzc+5QYvBXIKEoqlpBNVjDv1HL4W6vA4hbfqJOWoHHiGSIvjVr+lBciw78OqytXXrbLpCCsaa
0KmetEJntY4y7ydTlKTU+ePgVtwMWFiXE/mV/gP4RWe7JButB2XOogsIbLjJTfrE5VxYR4uKvx71
hV6laHrB1tRu++W9UHSV/KP4kb3nGKImoA2xd3xql4X4Oaj/2qLI3sf64ZdaVubcjHy12D2XTIfW
GuC3BbULTa7GiXDTKZDxbFCd8MNazAXeELfWMHnAtFDiMIuHfX39Xz77ibEz7Tt07OKfOktulc4N
Lhy/lwMfatLlD+g9m8CA4rM9pPmLLafaLjw10qX9P4UUmJHoFCQnrRAueCnQXXJUY5BI939zCAAB
iU+PbHt5sRkF6BbJ2hIDYJpPVk1v0Wmg1iELHkYaPHAh3rwHzulahjRAIojW/AeDa50BgsAYASOH
4e4lZP0NVhxRAiBbkbj53JeSZLcb7jYk0SA4oPSm2nSgigTDdkbUYkGxS0MFfWLXQc10MZn7zVIz
4ZSIxVKbs6cc7fegWTmENz45hzCNb5jSy6qHPMmQbyI2gx6jrbPKg7HLjVBPMRWHvsg0kPssxcbY
YPzM2suOaVnsO3UdN19p59DAxIo5grRSxgDzxEBKYzrjI+I+omXTsdfvOrNKq/9m35+i4vsBgWcj
7kTzY96RJmrkrZoaLFzge8G7lVvpwFEKBy3V2tlvBYJpBL0KfeJvdObnjnyZWKgSKnd9B2SyWC+2
jSvlK95uWfvHy2vmf2tACJrcFNkI7nStWgzuBs2UESlgacn3uGArOPoX4Rp0m2ZjqxdRDtAGMqaO
GerwP/UD7kmUknaF6/M6UQeXGoEBvJYiCHbJnm0f5oKKNVn874HYFeg5hBUGcNa5/gr9GvAscsvQ
jOSHYzJimefx19LZu0t55SUcPNzP2bT77d/DqqTyR8qcLMHfAACuGc6sZqSEagkeJdTVY2QM0dtj
lxg4kLLvExVvEEB92Sghjf+29m52TZLUznLdhPoi2ypS8XLjSNCO6pcLgYIZp+6ZDNhXW5UJm2HH
p+TogrFmXUboZ6UWDOIE8HGspwcEZss78IDjyUL1DtPRhQJTYeS+uENDHqfaQmrvrI1oIJ+XxJvj
WgdDL5yTc/cD87ZZcNk6unnesX+m00ZNv6hxUPFVQ5ABKu5PDMuJioLrckfISHJNNtaEmGUECDdK
yzzquX5p9d1fbYuik16yzZHGK4014slKx8JgJ6erC+aE+upxZ0xhgNq5PTqscHH6KekhCc6imE0f
DU+s1fOI5AU+OVGr6BLJ5HaaBaA2QywTyrePic8NaHTjub5WLx+In3tkRiTFQ53YmX4XViy17x8s
VXeILW9u9/tw2fZRG6L148Xqo7TeBYBGZneXXW8RQailef5ZHUbzsyW3iGcHZGDRqD5yBhWXSjuY
Gz+j/uMvy60vcNBwMfCRU5yBvq4OrDOS1NHzRniayXbpyX+Z2b3IRHHI3gS4DMxQBE2eoRccjckg
AqW4ifW7T0ZAG0DwQXpRYotP409VXoIisVd1pyAFDna/gSjtyzDVggKuUmwfJpAuhicVq/y/xGJQ
SikLNi4XPEIL6YWfEgZX24kVP4H1xO+b2fjVJwoiDSa3ktHJmruEiIu3pCWuS3h4shYJCNZ//VOp
qD5DJxOCwQo6/1h2WYOhZmrurRm+UzRne+FRPGF5wgR/yC4e0o+k+TzcXvKnP8815nE6sJDrDANv
4YHdr4hsGgnuVVd1hDHApYef2rWqM0aiVg2eglUF0Z09YNkvWjxird/bDphK34JvLeiFlbhFFNUQ
tfB48NiZ+q1JV6tLXIclUe29xYINWRipo070PhWaKF6onlhbckoXBYtine9npfV0K+2Hf2j1BvyA
rvMiCjPB/Qm8MSxT9KYtnzyYS6pktcn+sQMfUMGqURN8BeIgDB0aA2MavP4JLkMb9RHQLDknLuch
7+8l2329K73bRJH/BrVtblIig8zLmhKrpQVImP1TyCcn/9z7+K+a6loQ/vcuJc8UANdnw5wryKG8
srm9Xlx8A/stHRjZjB8VBTFp1E4yE4Gd/kyb6sKkuX+KLCsiYGZbO2OfB/XVEqwF92qZvvqOdq24
siPGB0PZfOdNILNphgQPBvpqJS0cK6Ml45VaPmDThyCQ4FtZbLvvefx4rEOkcbWpD1I2XOLlBxT0
exOrHY0eofZi0M5+Ei/fl4uT8mYW8Tuzw7tw9z3D3xjhpjN5yH7pxwMZusp21fJOo9M+zQw9VBYC
41tfaitu/5k8TylAWY6gaBozfxkvAxOyeu0xsWyuUzDWYj9+Ncez1/Rc7qt6r6l5T5q7SIdqPmF2
C/1tjflIbaq/lwBI6N/vAQmBScve9XCmy0CznoaF2omRu4RgmcxiUhoCeC1y9C7eVpuNZAQwQ+Jy
ZJviDXlx3EMStWOJdkpdZLqkjosjGVlaT60klD6VBLsZjUkm+VfR2r6JkFadwvnON/Fc3IxbFD70
GWWThPFjX8A8Z4e2Dvps5pXfP4WABQprlkhNpD9ZuHDSJFQDpBNqrYS13GLxDab7g1Z4UPp70rPS
Z1YOIYvX745g4Ci+7lid0jYrBRwRzAzWf719DxYBxxokXbeCapfgCqh7GY0HryEs27Vzde+zGqN3
mt9lDHpAxnw/tPQS58v080GmAISYgx/G7aGrDcOJVDtuL/uxNXdKcZnuUAffaOEQ3rYXbTI7ISqQ
aU4Wav6/UjX/vlT0xl8cN2bhZrVaNmt7beLNZXC51RWt4neX8HthN1ln+IyF1z9z21vEF6QqMfW6
Qs/YYCJWq2RMhIG7v2p5d/HD0cAaLbmYe/vVIZCV4xb7NV3JFnMDkAeUHrhxL30l/px6WXfgnF7/
2L35mHzJHJTjmj5NuhZjMFwOpYTwieyFo8bSck2qzIhgumBmegiSf67zDDaJe6HTWrbVAm0Uj0DM
pqQH3qsSaszTFIpIpz9YmWhzVJdqd2BUMJ9BmjuR6LkHCdL4TLdrxI9cH50wl3rV/mdGK7VSxgmW
56gyQ8xAoD3+2lS+AsB0JSeWwCyvq58YvBJdRIzwDOyEcSKqrdAIerxGDyAYVumQhQcI0UOx3QCp
qvAhjXyTWJTREpgJcsMn4RM07XdM0ll2fxmF8y3pZkzwTBndq+3l5A4PHSOio+1f+6RQgJoIsBjl
LLGDYoYxGEMUmZZLu6SsYz+yxOg7Kdxz60eK/a0j7ABoatH8iYTx5LeXrY7nNYIhoZIw+AqQMxRQ
uO/Q9gXtmq5i38QPPU4F+jfe98JOfLQEe3Qja17YSuiQCxTNfCE3+qqMW12l3Y1dcpvOzghsjMkX
iUVl4glsjiffURt6d0CvbaneQzJRZBV52WFxhhuKA8UomXzk+cURITAYSsbhiMjX7vnb4z6rTGG+
OhHwv3RinpXSJFo+TxyRUyZBZNuiiPhH4SbiOaKpNMzKEkMe+wtZ2adsaRyqb/7C4MZR/0Mr0DXO
bJ3FwuSTqIDnLp74eoYCOLIecd62rj2jBH6WqS5Def4TpzuE9dwv/4E/jtRIOUvv8zgaO3DWgFG0
hlsgScKWByphzu0LUJMfhvSFJwSKt2loiBSduEyatIuqGeM3Dy201d+aZ3aggI6DZDnR14IV/MXg
uK8BQ7JySubceLBmxYGs38L1JRevccO8EVjQyo1Z6OSsS13Zhu8E541N5LZDR3KzyfjTdBF2e0E0
Pkg5Yjg42DI0EgU3NR4lSnXpm8IyS7xYW36hICr72JzDt6pX1XqbDQlYenEJO+udmuB27NPXsctU
+WlN5P4aaoJJ4XCV5k7y4XpcwujCSjKX0DUWs2eaSLkV1DcpS4o8iwu5G9boX3mhP2tjre2uwNDs
YBkQIKFicm1erjNm8Z/IGbj05/aC+4G4j5/5pu/TSvGpGmiYWl/nv0LY+2Gps/emi1RDyW7KL7Lr
4MYWP+kObzSVEO9hCylGzhKVNGeXAgwykoVPCQ13g26z9py1zzXKf4EqXmWX5TpvRqwlQ65Ocvtp
HD5+uVikFAWO/TkJToE0lAZ8tHLMz5c6HxcfZuLQULJRddmiUAnR4OLo7Ua/SXL+lj3C385Dfaxq
UlIEVss8uReTr5VQF3Q7gtKIQLFlS5wGcChG4dEnnR+cehpacS02r9oiNVYAHUjJY+14NcNuOPuo
vrxerlFonmdvSuznXK2wjM06iVazko6asV04VdLjoySzuDRGJ5DP9NbK/Lv4s8cKyEB66N8vsuRl
x/cGbIh2CV2LRsvgzpfnfxzWS5MuShyTU37uFV6SlKapHxNzImuoeIgpFELkBKQgUAPsPjGQYbzl
0A7UvMv+vcVpGHYq6mG9//VxOVgut1wPRSoA45+wOmqmqwGsJlj1oY9IWkNxMTyddgzdSyBZhHmR
f3cQU/yCaWta923zxdJQslT2x6axVZJ2T7ofJ9rO1TbAI6bkJpbl++0rHBmynjEERDe8vmcZ3Eqi
GJOZ8/oAuPncEo+AiJPodLB4X+uoOl/CMAgQ3gF2oDwBymUnMaH8DDZyMy3kkgPC+klrzAEueLZA
aI1UohRcUO4wQ++Y+ZrAqaL5IVDzDnPFfXEI50M6ypFCPj8CEwwq8GQzBsMBHAD1zNec+chJzMLr
6UYx3Y11tsZIHC/ybp/c8B3fC2qFM82oJeaMFVTxhPuEzpUM2/VMphUb1NDpoFDha0dAn60w5Qoj
I/Fm8lreYtWvslp5z5SpmpNRTEazaL9Nf3n5Q3oVQWD/gAU4U/BW6pf08YCRiUJ1csqXxrBwuMm4
VfyV+U6x3oRgZb2xKXKAtTbRDXtnA0AwRn7jiOsFLsUiJaLUNSvv8iGAxI1If81VAIISTJlAGsJ3
9R0eEhc78egSsRFaCFdP9Pvl5ha7JAro618h9xRuGn7UeRBDDSQpFX4hHQ6Pv+hPDft1mAcXEzXa
ok/21ODQO+IWwq23OSxV3KPP53C53vmpvcBJwRsEWwBA4/Y0svKvVwBFwywJMjmvMvJ0HnqCyEhT
Pt38/KgSda64uNIgQieuR3KGMdHurPxmYXMqWATFaSrvjJYtJtNCYcIECoRaXJF1Lqo0KSQ9GU8o
fHdlf+YFasFe5gDJvi1gxFybj+TkxkBKWsWnclBeTSyCQG2LkI39K123I/cH53zoh9MijQdo4Srn
3fPXAXG4fvUfZA7TmqGKj3yjuWuNjPUAfR+tXF6ondZvTq11fKLnhp2ODRjrBAjbh5/ufg+Izngt
XzWjo7G5z5T66yRyc7B80HjiwJSrLQRQG8cGNa69GwnzYAQN08/Ha3Y+KBLP1Q88e6rzzy47bAmN
mqOI5Igc4NBFlqzbBWEc5M6AAhe669JI+AxA87DHo9gwl0Cv+cbDl7FdIFsfgudAc4uzBWkOhNAB
MfeqT0sYk6VXTmCyY4taNwV+j81DpMpHjjjvZu2fe2dvfhyNX31TCGSUW7p/u57Hm5RWr5PxhXc+
sWHc+5LQnVnwybchMwzSm6oFeQcoXBH/3xylwUIwncbVsEvk8jLJ8OkaCIFYhGk5CFqnaf7ct8mk
u5UVddY3e91O7LV6ZR0AlMeVfA0Qo35ghsw9cA+Y2OSdkwYhjqI92wF+ncr+9RiACweZNHNBw9aP
WVtgA/po2zH0XobGJrQgP5Ne/ZwHlDUxDarw1eveJ8RrTalYgiyNyqsTGNiPb9W2QbAfxFgDgMUg
0Wnx/uzPTIzRYi8K9vm89hPIx8zPajYU7IstD0xQB/JPYpGhnKRU/y4Zwq2B6x0nJ7jvB8pYbdye
qmiRMZ/Iq+U61BCxC5/gDLNoui+AXNUb9nnR32PBG0I6WutzxnkYk3ItLNj69TXWzJwb9MakaBf2
mYm6d0H16z0uBWXnaVm5m3Lf4iTP0lQaYF0qPRms6ytrw9QDo/i9oqRvGivJmutPqB4qF7n9ra0H
lKfwlNcIybgw/MtCCq4iCf9fOXtY2yxQ1c1f2WHAkztp6VHK5OeNjapyCLjIeYaEL7P610uaGDCD
Cujr4QT6DA0Zf7Npvk1Po8+pLzcK9bU81pUFhArT0vQe8xwVMJ6G03qU6W8MAqJnF/fHngF9nz9I
yFalte4S6l4tPkmt+7+xbl1eJ4lvdLP32AKTwPjcfzp7ipcJYgmOIu2kBhJKvPlc70K4xVSTifi9
ipNiK8B1zVBfvl0Bis2/bmC59rN3O1DJdOoDy/8N/9+doW4dVsY3xZZ5u0pw1fn9KhP+p7yBfoDr
K1gHnfd9YS+d4kVJY4YCpkdngMzyAZgpsMexmnj5YAbYFwRqwg6fmrkaPaO88V2vky61sA1teG7Y
oeS/vE1ou5u9ssP6sa8LCtjkrAa9hKQXCupH33zOgNQnGTbvn0AYE29qLwbjnBlClxRhe8UA03KH
qcVqeLApZicSrjVPhPvp13gxsA8Lf5q5ylFI/lW4vVV18XT47I+dhf9900FHQhzDfiK1q8qM2Y5o
yT3Yu0/U5A0MOF88OhTqAeW54o9UYfrKQkEB2Su4oJxoscL4IHk/0Qi2IqeRPCEa/PWzduRAtBHy
Rsv7mLj7d6rPUdDEdYUhvTJ1RMNTCZCyB2icAfA+tJyfYH/aq1la1TfDNhM4x6lwJVpqitbcqz7H
ry5ElO8FIWB72KPTYTirhZzC3dVSEKdHscM4NmSZCGd2hFGWwRgxDKl5SREN1C2P3R6RFB31yFXT
w/TLYd07fjLQUO1QkqCllq6kWECoJzi5YzYxXrlNJ03bh5kLLz0/r+iiRMpbRVRgvz+U73e9N4tI
t6CgWa9ZgtUXsXtXj/RljDkhG1oIxs0Wopt2Pe/KaNiRivhs8VlslkfwP23nxqK4czW0aWZXszfx
gzP0T9B/qav0eIymTZuZoPjwW6cnXrE5um+MHaZ7Jk0y1w6/frvOkBwfOuWIjK8Lb/kUqfc7IG0h
pt+IC/k0ytdN1KZCJVeN1LU8AuJ8QBea/iQeTT9YWP8AdKpqgm/ItVKpZyhj7gFSeudpis4+cHpf
S21i7S73FPKyDVlGlGFq2DlXSs4GoGP+atay6VMgW9x/7S7criL+4Xv2FFKqaKPa+2alByNglCSp
vJei28AP6ePFP1Mac43c2bnzGHj8eVRC4DYgUfN3C4xU8piAPWjpiCETFaWtARjt3EGeSwiNAQ6Q
0cz1JumC3ZVIPaOC+4zBe6lwS4VvF2y/369+hnerYIza6Gf+DxoVHiZD+HHoTtYTilyY1hKnmHdM
ycTMbO0eArHzhPcAIo4fmP/xOEjhog7iXtr1jyOqOX2jGkxy0I98Mv5NUbAQOnDe4mnbyElBT2dp
tmzo6UcAA+Ct7sWbX5zh4WZFPVcfAjzs+RRfV1VEHgd8BlFAOJUmXSSrW9e0DFyyoqdVpGbyvEif
OM0KjOD6ehBB6gvoE47/E0K2tZKqwQ49CWnXUSfMRZI6NiUltEoopG+CFVWQv2tQrVMZsum3TSeN
9QWwVofEWdSXZzjRy8dfHF0L0x/nzx71pLjkTJ2BMEH10fNTR55lTdOfxWjwN2a9mXMotN5sODUw
I27Yy8n7plxPx5TCNlIzqgEsAANhMWu9AWhdyUZf0JJBwWa4cfHN8S/X9UE4WCMU4b/RFMe9NKq1
DnMkj2rRPPx4QprLKVkvxf0AMlLmOrhGdew6vlTYSc+1ZtQOQtsvdalo2Dk93kw1tgclfsmP4t2h
16dRSCZL9ibBYJJB3Cmk/n6I3lqIkEd7S04x2ZdYNPewN45ntYZVxmGktmdFdK71lGQzldaFp498
Ln64hlT6X9hbiDKcXnd8dS4DtwORPvAzgKpei9r30L/uUrAvZ3Fzi889uM7WfYHS4skkuA6WpRTj
Jusd9Azw374pAD3mMzzdmQdprx6tOf5Op128jRP49MxPAXlmyAUxRMaKr16Kwa6oXsm0IEfsNEZE
jhMPWf9BRA7xsUPkRLTSyp2M2U+zJNViKmJiH3m77zY35WuNtXdp+QSgn+O2yorObPA/ISDzzw4V
NPAbk+pFZcwlzLPJoV4jvoMD2L+5sdW2iBOpW34ND0u4u4G2HAOiyvjdZmlzHo70FY59ls0uMJZR
NPcjXiVduLPoHPy1bqAx3jVyu97OEcGiKbRlAeZz0dS74qBZC458alu7bfWqqICYHRpd6eMncxtU
mbZ7sRqsCCyh7tu3eLzAOofsC5ibz4H1Gd9TogRLDP1oSEn0+KcrUC5GiSP0K5P33mXxam0kAjgV
tJZm3ogEeZ+71Vcepzy+hBKeyK1IEBnHurZcZvj/RoG5EinDzBXUOQiX+28sDXguUqE8eh3iJOxQ
naQfER+rinNxb9qgtnKB2Jy3LQ2g7RP8qYdBslfo+uVCIc5UIr62fvM3r696h4sb0Cjqh0nmiXzd
c2MHfeXxm86v26YhRaA30119YpCWeYhlq9rMa9nWW2wPfJbZuVBGRtUl1TNOUA7gilMsMd+JqZDS
AhM49CJYJ5VGq3LO2uLhr5Ji7fnQ2K5prGzFQTlnf7U/lGv23TODSC6aKQhiq8GkV0/rfrpfn6dF
NCD435jxc/xxXFIQiguWAAvhcb/n8y/vsoGMXk65HZfZKk4NuNJ9L9RoL1TLR5dIoRYl8YC1iChf
EwA4/12Djdp3gNdwaXI9ZfD+Raz/iHYBUH3yht0/WhBbpE40KA7JlbYG7ySAYLg3NZwn0l8YqXX2
x4yIonYyHN61shveo+xPBy49bN69Cuz9hPK4Qj3MRL21uxCDQUHIbhnLFK6XbWwogqJxVoYjkAaj
UDjgLC7POjwyrV81AZwqutWYH00id+mHxME4GvWD+R0Pjhikoo9aM5ebGxHtw3e0HgpN7igjhQ7W
rzQQ6nJs95zVVQSZghZWSnuT3k4SQy/CESOgfvZPKO68dlSHz9wD6MLfER4E3+DukjRPr6Ex7rBz
GKRQ36Rfs1uwEAivhuvPiyUvLO1r+gtJ6ilSswVVvhdVrolt8iZchaRmKhpeEbiFIRIbDMdCnfDi
E7hJtpSDPXTD4zlfPOBfAIqiK0YJtG6CpELNSweGIUegFpaocyO7Nh2Sg+AqfZGWv+6hBxYPnmZ0
LyGy8qZrM/0F/6uhEo38psxz1qQW4/JMPqoKp6N5l+YT6ZttdAnGMmNm/Y8M8L/atuoiaHyzUTQk
FDf31H6PuYKJgWqgZMLXWtdyvUVXYxh0aLtL3j6f9yihwrCVEyTGEhe0H2UlXzXry+EidYI9lo76
/X3hKbNQpNdZZoMvkoudVP85us2iFXQbDHzh2fkjwLWQ9+y/q2lSkoII6KYobAYGJN8mG4ADXTXi
CDCm20dzfek7rA3obK3pYB0Wp/hh5n5Q/l5R4ZdAcAVEjcUfQxQBrysZC3vPWPBmwsPGHX4gHmcj
56OJYGfkmKLLIJ9z1Uzj9kgXezOQUeiTWJBOPbeRLrJLr04XoHPSnqaCKCvlMxRCr5XC0GcdHfuA
va2yLg9KaOZqNgOuKC6gBKoGtefMqkiE7NuWbbjo0szy5yuPGkSUkZueYZdTvNARB7koyX7kvrD/
ASVtTh182OHoQkkQnCFw/98KuieFE1CPaOqmL5I4ce6vg+z9lPzXNeJ7EzlWirKtx3wi5UpB1vTS
1TcjBrPUwZw5EwGcWUdqAGQTjZ+5IwuFdpjf0TTiegk2w4njTVhMxwgjlLVQk3dq9gZRatFEZaJq
r74f9/jip2JpnOOy5E3YdQY1qYEDhvZDO62EIxmMsQEvNFOLIoGqZpkWmZ8iwJpk5/LanJQ1oM94
VyaKbBPFuUAl7fWCEe5PTR5LkANAEnaDTlB0+tVzJ+WUlBHeI8U1YcIHoSIymSkcquojJGOglmJD
QkRJOXm9Z6Io9gpRRA7xXZUS9QRcImS+Mp1HSkb1htO8cMVeNi4yhdqP0Z7F0sWbhgBErSLj1uoa
5cZP3y0qiMN6uijoBVQseIjbB/FtZtUX1xiuqGgKiSHQxwTXGSejU6GxZSknKvq5DPMWiRforApM
x+diP47RjC1l11a+003oWeKFR+8Mz8G3yKxGeYe5iKLRhn9eaZ5rFu+SDWQqwwLuqvsOdYy+GIFa
6GnrnO+XM5c0dw2EBeWJ3+8aetyaxvquqcLbIRnMsGC05WKLB5LT85y5EjhFP6prfNCg9QteqH4A
uw/Lx32J0+95iPG916GZuscvxr6IjNAT4n0sVjwlaiKeN9SpnDOSig0v1CrYK+1ipv+3l1J61qiM
a4x25XEvFGsdvpTv+GZi17iTjwDJCi1zUOM44eOP7bjNIavNX2tgxTf9MYOt3pK5rYLaMoD4Z4fz
dit5hyHuOCcbWhz2D7M/Jk0na3Ff54NU5kS4qKij4iWW/d4AyLxEjfNrmRV/8Fts3ZIX9+8OPMgY
pBNf3tr27bRxGQ6xOQxERapLSmHNtlQd1gjj1ip3mdjrjODnheqzGq9dUJ2S1R+tYka7LDNnKlll
bFQVusRUOfIsnL/nvCzaPaqlXjMnaxIapHraPgeXY0pqupSWu6icWkp8X9nVbC6iwJnMW8EMR1Sg
RxOM2RTNmcijocKZL/15eNWAfkpE+IOG+GeOhP6mmO7YQiHxht/c/1/uIC7F55/swsZsv/2a753P
OzKxc7lRjBBrUQ8JWDK8HbXg6U+gPvJI/K3p9q9WgTa0lVR/I4RzNz6J2/+qHcwLoAMk0/PfhWKk
0qx+pcdDxlY//EV2+CXiFtxK6Gxsh3b/F/sv2yk5bBaLfYbRObcotWDF4Bl9Q/NfN2qyRYP09y19
V6VLbybYjBK/0Jgcj3xpFDrB1qjs2ddEK2GNUfq2Zb6eVIIVuz+xveJlGM3xneIBKSP7X4h6Zn9g
hj6nqp+REQDQLA+VyBz1IbIhuhy47D9UitKW4fSh88vqSNmYH9erVW0O1G7V3+WfasK/9+mxyRqG
DdPSefF1ryJfAPKZSd3SvQqjAR43ham4ddoC2Z/GObZjc0Jq7Z+PTjMmc2A+59mxiYU/f8ADsRap
2PP0L7thgpM6iHzDhsIFbt8DrUS9Dga8h7PSS20t+vlEzXjp/JYCS/h5TySKrdS1eFDhXclqJ0gU
GRFpHEwu6WLXdB1yVMisn2hMu5PzzSUq79Vf5iNzRAtOlJlzICyFk6eh/3/MisnD2HCygk+atUAO
8MH5cs3XpfvP70W+qea+U1A+F7/rv+u9LUdjTXfAKJ00DOK4bkCOPDDPaf8ELTmPaWgzhRy6z/G6
H5N20SgHZ86x20lndS4QtKFTIjuUJKRl1HAI0lFTxNl+oNlQ2WO3QIkZvuAsN5yK05UC73bII6mY
MXXNM2G1WA9pwIP9QDa40KOeicT1MFBn9VpJHOLmzR9d+T8ipR5x0e2ajXSLiROFVda7ZxaHBkHP
4JAB5lECu8Nz3+xPSMclktIgmTH3BBuwfGWLbgbVXWWTkzNOIsbxsNJev6UWUOCE9GxxfL/7aObC
cBG4jFNthlyXj4XLRxDwQah+AoSL3QsW3vOOiLzNDQOreoDIRfqvyfu8h2O7+QLD1+WBfWdTQDoF
Jdav2RFdNa1jWIukk3aRcEFKVkrsEhPWlqeUD4IkRsWmQg+f3z0FK9w4+PQxRn3ds49gvwxIoIpo
nwIYz0UWBVkBR/E6khm/C+eGIRONSwtw7LtCeq6zPbfCiAd6ng0VPzwWHFnT+5Ltn6p7OrWBmrWd
vsXsTJfntWqnnKnFwDBvYL//jFBpj3c8odO2UWzaGu7v56GYFFZqmLuBssT3ujrg7CsC9cxvWnxw
eWyqh/0vTY/WVZv3iSFp6ve+2OBvOoS17o9wKlXgxQ0zPpGZACZGCP5+HTV6IHutWQc0W1bS3l9J
e3CtSMF9xIvDMU2Vy6q2zLtn3aPbyJuJt2A6Si0k1t+9zILT/HjfgutYDsUcIwtp0ustRwzb8YxJ
8m/UFaHRLeRGXTK2twavQ0eCLbkQZz7UXVLhvJNanrLUenpS8pVR3a10neCANIiVLI+mzB1T+naV
AwpGkO9S1Aj/l1e9sdL5c8HTvNSokBZpHAqI2/7Kw4825Ei2Mr8CG2VD06udEy0d/QHLVKYCEBDW
0/0HY+aaiEtsqDxDh6/oDQOSEN67WlIM/aPYsENBke2RX3GNzb2nj/sJ2BrNxMXLfS/bFqX9U+wr
dZuv1IKRzN1oXZqUND5Rd4Oyn1e4KPO5Kcsl01+G6sUmlCVy7pHpcm/dV3hS1madTelZmLoRRyCO
pv/LGS7M0HG07muontawUZR0GFytHxM4Zf2zv2Oa4Vr5Y6IVWKACWpIfVOF5I/7K6vSw5sTVVqiS
rCzFPzsiCVR4fqRJ6YjWNPWUaR8nhuyHwUY+OnPbKtVgQ0uyJmG0ip4bUUKapCBE5R4N2BIADaD8
xsBmyx2oNqHSC8RIc+vTu+jJy1g+1A3wJOujNBYbDWLGzgk5of74Kh5JS5doy5aLSjW5T8wgDQNx
XoWl6YQLuS6C/iTzAU1cXYLSHIog3MNZNX3Ml4IRltZb+6ZVVBPtImMPwTSwk9nMEinJSpZLeAJC
XQbq/nKwMsezCnbbMIYZ4lO3gPrts1yK3HaDGiP5K5meFzqFl0f2YwKmEaasIVwmNtZhRUcLtw2H
IvP8Bv/F0fMdhH2m/1HDGHg6I2KQvfHjbrcESFuFmCmdmGaP74CIatq/wXYwwMJy/YAvPEIyZ8v2
5XfTys7DuqZ8FJagMp7oAzTs4Dsd96YYSd0Tq2UbsZpllPi6CbcvUfRA3OKVngrJW4QToH8DvGUr
c3BKBAMEENb1NLqGtlNUnr2WrDlkezAoq+31QxRgB+0+M5QnmPt/jik0BWr5m9haFifve04x7Z41
pfDRctBY4hNEDyBEPSzkWoCDkHDth1XrRc4N1Le+lK5f5NwA9VfjazSsRtiRkRaRRuCk3NFvFq/Z
Tw67logB0DtdQOWvx2Qsfm3MgD/7NX6CUGy4PsN1pLpMxOpSxpE5tEbN41JgwRzy6woyQvKiBKuv
AA879tklty7TGK6SEC0oK7KtHwUQBO2zxV2pUwlFrk7Oml/kB4D+i/S2+SaPDao5ieYZAmipKgUv
uqG1vFn+luiUbMu49bljRCIrUi9IKWgGeZP00/wc04FvZovsIFopXlANt8U2BAlw3EOsdX2VV+HZ
xwb3XC6tlCO4lrKAhH4zu16eD5L3UH4blLpxf+vQ9kMhL7mRckLJvv/t3LGZcuanirAl+10XBuJi
3L09zfzaNIDe2S+NjZ5ittyD1iDIH+D5nu2pKzOLnWUGKRVwTaKCCPBKOLfUhobtxul0bx7L2TGL
hrSVuEpON/oKZcS6AtTpETFBMokTtBwzPma8osIK7F7rj8VvgfIjj8WTQ243SH8lvFGifHsSDq0R
ZjhohNELPWk3qcWXhCrVU8KxDFEDHr8gGeS7tp0aalg30gllzP/NK532uWNsX7OK5xbr+cgpM1f1
jJjmgG++qacHrU1euNPZ48+f0IKtQrx7WSV0pNEZzz+n2ENe/RWzRdbYnHpxDsKlT/YX3FqLaMB2
WRIdo5r+3Hpc9X1AOv1BdE8Ov65EzxZn0/+OTaUjmFqcNl/bBcoElV2Z5rHS2FLs9ReXaLhgypfb
lUjKnqa/gbhuARUCILE1bX8r1lYS1+tWhm6Hig0aT9wNIkQJLWiPmlM5evsNg1DDK02KZvciJZsx
7yy9gRVc6hrY00zWTRSrjZA0o+avjpilCOiO6g4O9c3VpXXZESQ/QoK5+UkILqOTYuzkNnr/O3ze
N82nsHamgK1UCFDrLDqmFmuFQNu0qnDxIDGqazR5TF+GdqkxqSjv8WEf32fIFbncoHXBj1erAlHL
NUVMlh6zzzNCkYXcvRNG88SblhakaGz1HqNPVzE16lqS9+2SwuhAXsFFQqSR7FfTUnizCD7D0+ir
ZWVzvIc2n59IRfwHSXIDOxSGRAhlb3x2/6eJ7hcTSGE0KWEvDG9cEze3iwvi373XvMSr6PrVYH21
TV9pjBzdYMMmnMcSZfRBRX1+YYtSgTQEffoWliYqfY3rK9BrsKWJ1uPYX5hlzb08aqXly76gzIEl
0T45UVx9r6J6ThSxr4jCplkirNqZhBVAsoyAojIwLqKHn8NhkMJT/qUNnHsZkT5Pdze9/mymzKSm
vYK/kXw15ZH0+x6lOZ8lLXXicmwpuyu9aaax145Bas3XHaUjy69H5Z/Z1ky5ulSD2gUYgWoQ58ip
XSq4PMhqJPBWOfyQR2JnWu3ZHoCQHE1uVO6W/5keozhpvrRE9ki6Bs65RoZJbNeOx4iQNQChSKOM
9Thdf//HCv7IJiXAfNo59JB0XcTVCZ96Y+rs73GnlpLnYALuAoT6q1Rz3qqW3sZjBWJ5o+Kew9vk
7wh+yOihEy+24rjIBhZS4UYC5A/9DJ5IKLPm8WbjUaA3vRVcYPbxMttJwjVe6lBhnyro99u655aL
z8O9l/LWN9Twnv3zC4swd5PgGsxeYtZKGOrikGl6UyYbn/qDUI5B/kF/4uEBUtUYKD2BqEVKSAOU
pj63XvsqEKQ4zIHr+KXYBsCnQIMfSJ5KrhIq280MMyl5fah/9Um3n3tfmD3B6ujgu7y95w1IKkdT
a0GETGZSyqme94QNhi24iOX4sED8/YCxu9/sw/HtDBkOLYSeEdQsG3d6zGnyU+ykaXHAQfDljZFk
hhom3oiaMssFAXIgo7UaaaQK0vdM0Uq5x+zD0QusEbyIEceCBJYN4c5+RhHLGW0Se8J/gX2ROGeb
bZ5v84AeYh+J6LFZW/A5BZAvJ6niJgxG3zSznQeBzYWr3Q1cEJ9UDooP2q11o34FDIOITs8Z78c7
nzk5pjH9wVgGzubr0GCTGHudmlBCYhfsPN/h9Q5h3xrIJqtS7ORvsXsVFriUQcJy/23UpG36OAfl
mHnLzyvI3CozGrT57MqQtqLSR4ONtEBpIpWIpHqR/S6bCw7vS0coNkYLI0/r6Iw+vL7taLuVTHJQ
OiylyxiBKtp6Bx7+6Rb9VKkn7OSBgX5wv0DPdivFnXw+6U8uc9OUHLmv7m+QgWJTX+Q4vBV71ZNm
hWA9+ASimY9j0SekZoFQi7+iMBolOO1YdFI6U2Vwsf1dv6OdwnK0Vu/4N+uA6dStlxZgTy60KV0Z
GmyL3oFzg8osNAjkXfePJD780HjJNaH1dzWcUr0qBW21IBhJQPcj0MpdnpfPNsiCpHai+wvDelYC
xo9jh2X5O/58PKhRPvKYR0lP+vtIpT/IbJatvXo4u/e9Dm0dw5K/38cFT14gQ5Flk/4mYxzPa3ZO
D6cw9bF9XzCi7pEND9omsP9VpE/xaryTFbeq4QcNE2KJuiW1GRjPv771TABSkSQF7HxrMivFJXtc
wpYALy7Q6Ey6lLN+iKYyZpYIL6AdObaoHfeVq5a+ColSCs/OnRhZZ+nu+0zJ+J6nyYNS6Du+RWzl
R0otbVLsOvXl82QNIXSayUVjoFWEr7Z2omXASfc6v7dV8WmECueD/MqZS2RPZ2nhIwO1scibpAS4
49dKW5HRMRU0NztNLFgkdcdRrzejLqIy4TE18IVaficaPcpb6TS8CTXD7t7Isyw2GDjC/XOVkccK
7rTvrjaJphk7m42wjmLpK07lv9X6jacVwSuCx+bE4ata2/fE1ttIjH3lyu50BjVGYXA+XJHKie3x
fMXVqFYAAPXQVHfvqC352e5xZy7OD3rZ14xBAa+Zy/cnQhJ5GLCAiui8bt2Q18Xh8Xq7UjL3mM8G
ObD/9uO0DXr4OZrmB0k33PKfUW+YVpgioE7oY2VSx2iVBtBghBguacHVfGheIsughvRrhBj6N4kB
wU4tTNNqwBg/T7Kcgyr/Y6rEkoSvWefMAtAuQ4dMCGmDKHLVqs2nnp1tWZ3/Rs8lncWnUf5zSafK
NsNFSzBjaSMABK50XTHgi7nGESPTS9WwWWO3oieejzGyoxSBYCN3E9Nqfix+QK7HQS4i/daz28f8
1XCn057USke5hl6Od3MX784RSIvH7jQgwRdLdxgVlHUnwhXDJdv46SecIBr41IEC1cvDg5fUwyKl
WOZ0q4CRzpn7FqyBISrF3C2G5lx5YnnyANvMITBF9Tu6RUPW/uYWWKUs6jk5pxIqDW64d8AzbTDl
vJq8KYe+zpcQp26fHZqZlwIwlGzuBuE4Enma85gVLvuFSzgqtK0/7DXK94H/CBLVGT3OCToqtKLR
45RHqFTQPuCicE9Y36ezRttGHIKkSxW6YXUBCxDo22DfueBO1xA6i8bQjP96cxQXwClqy554SoRW
3cMJZXzLspYWBR4WBMkRzB7A5fdF5TPqejviO4E5+MbLv+XQ0AVC1ethnqqDQxwyT0x2DE+HxCAv
4d+K1J4g0DbR0+D0LaK6908z3d/2w2uww9GZv5veRY26Mv+Z33+V7jAOFVb9wG5KmxHTkguZC3Jj
W4dVhjCoIPtL8VjliwV1CIKxZKbDrdBO3OGDHETeiUuYlyNt0lvW2Eu3/J796gKCjeGGNvIUVYby
lDGnFth8eUrK1H1u2RVJstxerhLKtrTkTkspFZojGz+IoU1NZHAXq1emofr+CZc0RyfTXaOg1Bu3
v2L40+95UXra0MOcKrkQh8hL6un38HZc0k6BRpLBP3IFzBmclpEElJ8hIu933mL+SkwtaUhw7BfP
D2+y9vYraqEVoKbWJTkkE7TAs8fvFxysZht0JxXvUZgamjYXz/oO7RmlMpmSNnD/Pu4f+6aGO9r5
I8bVuDyk/eC/uvUiuYW24/Wyb+tGEVhByTpqWHyhru8/Zf2/5Yu6Y4y+yalFM1qf3Yc7vD5Qzvkb
oaHjlRURDHiUveEX8Fg3lDxGbea7eR2Cg7d3unW/RrV61UeYjziJ2Wzq2GWzy3hrwOo4d8A1zGXl
7wSa8zgJjt3lnwEDqDuDlKHJuYp1fH8JEfd7epYSDCvn9d58IZQzllo962QanLmFGahb+qNVQsFs
ET62erm8g0V1FhlZMPxAqqScSFYtUwkLKo9BbVoAw65sCLIibi7Nf21WUrg6lQpAYLxBo5MG6G3I
k5+NRLGwqRXlaYd7DwDdEYKDtkE82MZPye/AVqIAuc5fwvIqBgS+ip7a4Z7VjH4yDrS5VXsqBSZS
O632yMWtBAMQ2ScRdMEfdd4mAm73bgApZXmPxxy7US72fFWA5tNF/n1zlW4HCfttbDK+iul/d1kr
lqzCVAi87vUk+28KXU5gjG8pDP3gwhxq/HKszi3tUmbKUzaG/Y8M9m4QLPnZSXx0Xo6REXHInrcb
FoBqydX77cp2/I/RKEfZVWRVC1gWIvB8Z3Qe6GsljI2vx0ZLNBvzxyYKWSyOSx2JBnLq0qnbPYJc
1iry29Ldd4cvXiNvXAUgHrbz8jW6ego6R6aLTUEBHcqZRW4CwC3sRRtZCa2BoLcWbyr6iqilnQY0
/s39jjL03wUnBCtm5znUVu9XDmsxGLJr8x0xTrx0H7EiYWy7Cv5lzdS7F/WWSbFu2h4qpR7/dWwL
CjEUnAZIL70q/NI566hQ1M2WvOX6e/n3K1V37Z/hkruGkI9Y9Z9A43Nj6zMsSG4rh6cKD570t5bh
GzMrTWiQeTulflTg8xFEHVhUQkZaDj9H6DeIRbQT1427z8FN+T0D8n8u3RR41pnZNx6e503ZcPvt
vGcgQrK8uP8UTENKUalHJqcA2IU9/XUsiYzjKh3hAKUdQ0eY9wJgUo66MEGceeVfYnuhcbOUKhdx
aDIfktSEP6uyBbvMrfym5goC1QAv+9tjKmSKV38vNuV2zkdUiFC0tXaR3onY/cplKiLcPS5DSKjL
GkyGGXGfd6KO6idgAcMWu9SlGUe2fCutnu7YlF/toK61lI8bL9o+Pv3M1Ilv9R0u6iKebagavBEF
qIKGiyPTUTUsBr/mO5ccerxWhBUG0vaZug/Xr8CZ8RHA1HLORDvJ1xyMM3jlhXx5q2/txpoKDs/Z
eeckU+NneH9Bt2X0qJU91OiODUsBGxAjcEn2s4vHPQgKjrlCIz/d03MJ0CmTZQpjR1/cnl4VgDiK
tHkR4ITnbz1RI98OlIXM8syU8+P21SJX/BSIFm5MhDl/XLkllxZ4bOV2XaF50TSGNyRknHe5ZFr1
2D50pAnGl1rjP7HNzJXOVNZDufDpfK7LX71HdC5ombpDyyGxu5j2uzeVnRj10RZp0AwK3mnHW7sE
XClRfifTxRnq0meGrVzIbjAG7mXTU7VMs9kwjovTp4Rzra7lgSFMAWZKiDbArF6Mb7JOe2m8+w9l
w6y4fO+DE41UzqTPwQLFQ83euJB8LUXKeNsjZHlShqp1ZINUPxo4QuxQbX7BzBJBmuhMItipJ6wt
yUxhDhcdfu6ucMHWPic2evX3ciUtjNQU3dj/u+7YP/L1TSkwRZljYnka8cnuRhFnvVvYMTwL2H5S
wtrlLVA9foQ7xN64QAP6lMVuTbwCBunVDZNshh2+HmEt3AydjCFBNYSEPMXD1cYKqU2k0WkR+AaO
E3GP0Y+Nf0MFKqFCwrqvBJjEFFqK8f9GJ/Y7gUntd19YTlAut88H2lXH2v+JtUAbjy1k7EA/5y7x
czdrpfzmS7C7FDj6s8uXyDKQTzwi9MNlEnPgGRU4KBFcoD+tNKI79gyuMASqAVrL45BC9sGGj3hO
sU4hyp6ryIVBSllLm7Cc5uoay7v8S6O9GyrVa3bIUb9zmxlH8uApr+MUVIoK0T8/fmR2E4XrFYmD
0Gv1hNGj+nqOPYCMqtyGeK3UcGnplFUHVq5Xg8VbW08IwR376ohjDi6lU4QRZjP18WAd8zS0hBV6
+qvxyTuHgAmqB/ysee4XxZubgUmpUa8Dh32J9sXwhcyKrgFz6jblnRQD589j17OdfZ+GzGQ+ySQz
5wAYoBEQ7LyKUU3CQBukkbljhTDByK1btKTIk5g1MK7Aj+YPTSgQAbYiJe/bhynjLZqgSWqWlLY5
oanu7ZAC5crpb2jU6uar+DeCpiOl+fkJ9lfQ8gTlffax7asRT6LLfjcR2a0bOf3nDZLFfUF86zq9
dCRcofZHbVU/b7bSLCwY6zhggNYfV66UtDGO+mro12GCx1+eqze7oeTrO+0pNncxMCbkklIiSe0U
mYnjxdxE3OWneJZW31kJMjp9Rf33o6Ntw/2UodLWIzZ58rgHSDIf/xKxoPTAoWT7LhprZpN7JQKq
p1uw/EqYDdH111gjXLqc63kZKVmlhzu2Yb0prJNIKVSyVc04zcOs/9K6ggEe7KgoTwTxp4DAGIzF
pUIIrgoMC4JqNvYGJ6jsEtkSTu3XGcIgE4xUYlJf4NsYtq2NCnOgooPZaTVrQ5a+HLpqFNYpykh/
fZAUdVYpEoOCHsTNR73sIpIVBM4AuNlZTvg/XPUJeGrrBTEk+VPgIINehm8sSQaukdYlVnm/onf6
PKfTfNImqo5t/RWYOO2I1jthMsP4UBrRo9ho5r1mVg6eFrQYzIiVs7V1B9g0RKdMoDh3cMSSkRPX
PUQr3qtjYPISEMjUk8keLyCNA80KwhfYWke+9mz/XS2DENUiiHEqJCnNbTQSCBS5Ghmf7REO2V8E
ESaBNPw1QoQb3MTx+3D8oLdU1nYzrKefLYbY6TDiK0gQrfS2lfG/k8Y79JmkwnIgt7+kt1gNBm8P
+2v8nksDKkvTUrSqLCy3d4jdFo2Nv19OVi/5PODpstwIqPKd/u9D4AhcxSRxoC+Wnh3QJIqLUS6G
STS6+6Bd8Pe1UITn7MVakfGYWi0Vk6NwetSw/UkD3VbzyoMmAhlUBkwTHSAe9Nj148F5CrCXGwHt
gGBOJl9R/4isJY+JgMm84c95YicX4YwRhSVVXKcl2voZ71Wcv2FdWE3mX91eGsv6rc8QANGio67O
FfgLN10leBU7GF9RT21hO04cf9MD3LI15w+iLdflYBmy5a7mDPoeCV+5C1gHyKBphBkCT3/jKed2
HzPFThU/7ZaKAHK94J8zcYo0PlEnHbqB1OAxaRHddaZZyat5vHnGDQCjkYKxDGuQZajF54ykUDMY
Cpr0aBjm1/v8H7NLiLAVYZE6+gnOQy0sAAvpWDiM8k5x/oc8owWgv/KvpXymTVZAJibTkKIKu5qs
JytztS4puzNnKDbr0utsMJ+wsbzWpVkleZ1VkAwDLCHcbIzOvTI6CkPAOmCpkdfwH0UQ5aqRGeam
e2WMlG11zeWmD9iinMZ7wRjcB2wYy4QWs3B0TEfDtG+gJozPLgAtad5/u8IiRI/hGa7HrgTGawmk
jPtqejPDDGro9kwBW8Abjv9I5Jswe+WGebIxbsuxc7OYXZONVZlpg4OnQgUxNxvFcQgY9iM6+qbk
XYysvyinKSQENpVGtwIuwREJ3/japP7q1iESRDsbRLIXRBMdAcx/UJXQii+yuhFvhZ41c+KodTnW
sbVDDp6HIa2ulz/FU9cVS73IAhQwA16P/vWzm1jgWS/t4qWaIvkCQ15b1lScXsKhu3Ec/PwBvtw8
w+knNeMt8hw3fRjTqMB4Liro6Q2v7aFDxe5u9rdTkzzFQdiJvCL281Afw7xbEGZbBuYs1nv3CYjT
lE+B/C2yPrkH8z6B9LB56Fx2gTaDClFuXapeBXv+UBxnsMkdyiKgvmnvhq5n/Y4FIOBgsGGuVnKk
vXBDyibp5oUZ4LPJyoPvH9hIIibqgusigx6tZ9LhkhXQoh1R6IgmBiiSakmuFe/nb490IXdlB9r7
t7mEuNGs+ZmzeDKSOoiBI5HJ7u6VSL+5VjXwWp+NwMmiNG9hHqttgsRbAfLbUHJ4kqRB1K93Y35c
lfUdNLyaRgJk7mGaQ+Bq1p/ickX2JIFN6Zds1FrpitdnRNxvbIVug1LOKO/7eS9PZaC/KZ7wpuPE
ulXnsi3yv/WydYXHrslBANwCVqe5E1BRKg8/rMk+FyiYGdVLIKwG5hwAUNFgOQfZ63Udafruq38J
RyRjVwupj2g1Q0ms3Pd6ZQQmPjKfdGigXnlHNdIGzEa8sf/3ISR+gxFoYst66f1CAbDtdxrJS5cX
crMSJIvBPHTzVLN8cCSfj8JnTNdkKbL3/lvrxowgJDJQA64tD7cmCjQw9sD6XXjNPEkf3f1mFd28
LikGJxfTOZDuW6Qfv92IBpXvjtvzG0dVaOh53nhKgzsJjs1slVHEw6RISTdasCg4FdlSc/Mv/D8W
pFVr6AeaWkrPJN76SAGwBAnsus1q9V8zPBcZWRujaVXN7KW9fGAFwFCYp1DMu8YDqw4ACURnYKaw
G74G12Z0p52+LHuLkRc7DIjhcg5ti3pv2ZTJ3+Iq1uamdYctw2hWBtMJd6lqfPYbRIsWCGPM8CAG
H8ZoSdByI6z67/bZfjqjESE9U7lfnS9Uk+sGjZOLf0ff0cdDXCLDSXrjxpkbVWUDGlNePiLUqGZ3
huWSJdJNhrvMTGOWqT+JjNYBlI9qYFGab/Ig2zSlnyJstrISi7PYSOVYjBiiYTd4UuSR8aEAuAsY
LjASpH0ul3HaRYIY45LVrsllRgsoNtes2Xe9ynK+TZmU3hXD7tFuGEDjWvMl0bM7l5ivVTNMDkvj
IJ60HcQc5+0EsNFYXCUFcvHbBoQM24pH7OS+801NK++tTCF8cKwDft0x1r/GlO2I/zUSzvfWLzjR
lcFMumI2FwNprLticKPuAzw/oHeusMHrhi3HXa5IC2gcxe7tNoHqrqsi5qdMS/rNFLAywNZesomo
UApwCUulz5IY3SJe+ZYEAOeA7jkT5iy7362JfjP7cA+Z/uX6YzJQBXRMW7w6RTTno489jAJSpCHn
QeJVLj9CczEXy+yGsRwPHU1vbG8I1a3KlShiGHfC9dXDGWvGT/WAlah9Hkqq5i1WDKIdhvuqkrgA
+njWgB5FNLkk9sI5q6GA2QoZWlq0B63eVubNq0doAfzBfy3bqT5jWu9WPiiLr+qZGZp6u6IQRXOD
45PEs5qHKgl55S0VSJKZB7gSyijl/1e4B0HgFMYKhqdBqjMA2zmqVDmgyo2VUmppIWxqHMpwYxj4
9p7Z8XBmD1F32zaaGARGdcDC3Pmo4aTFJaqhLsFEIRh6DkEVgvJnSVp3h45RSv4nFmfGIz0GosKq
LI/LKnqfheruqzROH6pf4ZWFJ3ckf+SiGH+1jtufsQ9YhA1TaZRPsWIm4Mauwuf8Rt1G+4S0G9kH
9MNABGseBtNmGBxR3UKFrkGIDrFx8Mb/vSRuFFTIWDpOi134xhMXYJ+19NXbxVgXKUyWNpH6g+87
D/GW3UHzTh3j6xAD7uqzsucK/Gv3cRxfWYl1ZVQk1doeZAONU8D1DHkSmnKOBMdPNNtpYNqx+Iiy
2xyvAgbL0BAZh3FYdETQdyohIe4dhVqMu/EpVua8nNoYgGx2C+HX0BMBFWeobGeE8lOOdwKD2zq5
yLrYKqbGXIgUuhA/+OoZNpOvjaBFfVH20lK0wGcqreZK+wpy/I02RgrtCUSscIXkxKFphZV4pXX9
8EbK4K00etGqyB7DzkGYVz4eKgHBwMSp+sslXr63PGuL7kGQ1kfBMJsYS9DKG5mBPTZHxIDSAzex
EkU7dmGa6yRBPwpAALWIbb+WPp+m87xnNCERJ9jlaUf8VxwrwA5sGu0Wz+QxHpgdA83Wf/17aFlq
UGkfSovUGCRYWYxGaiYSEP/mBsTVlmBq/BBaIf1tDaSlul6SmhcAwSnta+pZILVDJuT4o9knwes8
ClMgom977jgCCZhlCU3ZfQQhWjCbQMOrzD5CrKqxuMSUmhICDKJDKyqQqazdgx4e0qb7nqMuLFzs
qNX8ZgQxirVMBE3OM+C3uQ3ZFBpLG1dfTR0tbN/PaRAg2Twe/O8UhavGDnl1ECE2w0b3VPg8CV4j
bHayVcDIYXIfbvbt0mpfAAhuuzcO6DvnNJVS5DeMojsDK+ePOb/1JX3xAusKaScAfJmhTkbM4biE
36pnlpkfJO4yxJWSH+Lp2QBVPcI3IEPw4/0s4Am0ECzHrK/W7ij5GUwdlr5jDOuVBTy6Nlutd1BP
Pb1qWyii84qZKby/65Xl1/vOjpgHG7L+gIjKCEK/EkbEaMyqPhfHZPHKXM8w2Mea4RCaxXM+VKhi
gc3/EaPo35UAYTUqLJVuzgMtrSPLQZzjmOJLmGmAvMlupPi2hULSiWxXV7P5hVP1kZD5jqrf5opX
0wCUVVLxkoHdQfhhmVSdQt/3fm1bCWosSdJWT1GMFhxCF0ggQQ7KcyLSWYEwNpi3sP0dVwDIcCm0
2/vppMDwvnfZbo4kE64T7tGZk80kyXFPpCtvGjL2+Z2FoUSOo/91+x/KPnU+2DS0Ru1afZ0asA08
ME477I+ZVlLb94bR+1qfcUtx0zV/soKPjvSI3ockQMzrrM8B5JGWwN/yd45azkTgBP0a66ExPUEu
1WsyFtlCuCjHQU7u2i51/qgEEB+XpGZlzupeCM3+2RLGqc6lKCv3EXZ/N+GEYB3n7lKP+S0OHqiN
jYNSCySp8cIuB8A2EyPhIis926UvRkco1x++L5LIC+Q5eaYawQfbnNAim4rzrHeAjVXWwISYi5zP
jTVqvp7yzxwQNqrawCm9Itd8VoCPY8nfQsMoTuS6gPugDGgSe5j7ACZ3I1OfMLp3F/RTUT4H165f
vGjMGz4tSpcbIu2kcK4jF3lGcOH9Q+xlxZkJoSpv7dVFoCJhAq9bnB5hiScyP9I9A92N6K87/pLN
GeWtPJkIc/AMAGPJcxoNkYyDynndkkmOQpWomt3mZ/h25f1KpfGtMPOpvBRKpJnYUrVVIC+Vfz9j
kNvcLWx9Yi6IAC6Nrk1KUTe+6QTHT99QxmtZCeRLmIOvJb4cli2Xedxd/oI7okh7DrvroonIjHHO
pDg38StniH5N7V/M/Nzt9KUCcjpsZ8JnqBIApK7GaM/AV/xgCZfoiXuGkW+8raUyiVgzO2ziLtqh
dDgWpiXWyXtqPa4XHSqbtgiovVl1dX3E/IP8E3/cwAmjBwzs2URq0Ufbfl1rSjHzz8cQG7jWMuRz
55DIX6YN2QckQWq1TzMVpzu1C6SHat0YNvGnBqnr873+w6Q2MJqy8RalzX1AhrXjqDyW7qaEhaSd
RYR2bISW8wtiI7fPKjhM2Ho1/0MVG+ysAN3Mk543HWLT7nrk1vJNIOq5awYWB0i8hcR3WCIHuxbd
kT69s+txz3SfZsqcI0yP6rA/QXL6GdkIhMm2VF+7h6Oo8miuLTiPIIV3d5zxs7sDbXCSrBrlQFxy
WdOmWZwym/8rHT6NwDHttd3GNw5REN35mEBoBMLKbOe9yrkMmuB/6fqQuhz0K6aZrXJNkb/VgX5q
eEibZdThb7kjr/fP3JbUU79QiNYBtyCSQk9k/9IKCP1ICkhZs4O5nGrcgwpe28OJqcpirWxCPjqQ
lMz49BIoksDlB61CqcdfvZn4/JTrOXV5UFGZhvW5K0HZHvHTRccxubhmy6pToB6BAQdVg9pQ5rWD
pmES2suLE8P76xW4lBaJppwuW6FOad5C9rp7yaZllJ/JkkyDSFZL9wccmFRDRG+y4bFP/WVfTFfE
5aSZ5auLlLz/jfowIaR10g4to3+5H58omWOKQae9ZIDZNNwDg2ffMgjPdYZ+A2mJzaZmRFKe2kMN
99WRzg7UuADNEM05omTSsObuK4tamUaT78MqNaQ2LE10IKB1MdGtNequ7sOhN545e+hkMrDJR+tq
ZxjdO7oLfIXWKW9t+0UD0jU4bkhFNhaesOxYn5HYnCZ+7reZPWnNzBBt+FxTLjw4HeaOjVXwA95A
9zoFTgA8Pau8VAkpprqH9/7h4oX8QMftM3L31kZusLHCFBy4kqYmoIUFmu3wgNf5AzE4Y54oiXe0
l9iubStFNz0gIRCmSOv9dCoY/SFut7KRHSsMTDhI4r5etPrJNJ8UwbfdLQr1J8M4wlEqofzrP6iY
BI3D/SwLRX/gLDIPSpNzaqNcilL7xKFQxLlK1orM1ML13tIdA6PKoBRUrlkMr1yOTPmCBTLBKYJ0
3pzpGhJmAYtgaIOGlLAYfQrmof0mcD6fdHzXgMdHgJyz+nMZ6dm+tGVmBW/XkHPKAfDaRtuipQpU
bFJYJSgPB4/BL3i/Se9m7mW0RSNjWJHo+pD7rh+mbBFsAEAgskj7h7wxshologj6fNXkBQzdGM5A
YKg7PZHRmDGcCsI74fUHAY3QhofjOyFemicMeP0b8FjYxEUOWWnG4XBdjn/vw+zVIAlJ26ke7iMV
VAXt7UPdHVKR0wj0onaHJunzvTcX3sJn72AnNGcclUA6jRV2wiut36r9WI6JRI6o5+AFiYtMve5j
4NP94HP6XBETOSsrIUVZl6YAbTnKCswj2PwjWDsxmg40v1W5qvWld0b7l0PI1w1YrTOc9VfbMcGi
aRESM4vcHEZ4JsbTMebX2qgWKIEvzW+EItpnDVLWeH/KLFD+4E+axbmYSY9/sFF+c32mntLbx+Fk
9NGnaoI2cyXNYDl17r/N6Q674VWPQJEzKn9GLSmHYYpQcluWSpLYUEnoIPNtf3qThH1+Mh1yIocC
01qIqyzdpyhtB96niS0k0lteN/UlRVqZLZ0cmgzMAO/DYNBJEnaRM8z4DnRvGh7kBePmV0kIoXUJ
IFzpgPMKjJWnCjhNO96v6tlFh6zrLpcYlmsDM778t79L/Wgi0qGxhbXk9U1By6qJQ8YeqQUVmIVy
E6vd2Fou0jU5nojCx/4t8G9amsiQOT1DvtaJyIryOCIdD+JDPDiMGrdO42Yj93EoSH/oMqaHvpig
QhKG9zAhIMbiKo8Z9jRmwSqop5zAB/ief2PjwfG6U7TncKWo4M/vOL3b7juOpq2B1LzmXOnqnhs6
fP/JDurI93Novu29lnWbZUPKhSzLJhsWNpvdRxGlJ4auSR53fGhXzNJ4bS3F+tdWr1SkFr8yxhif
enoCfVXvRHF3KDKzN7hDqLk9NCQ+2iQu2bnBNuw6PhMJ4FbCdzg1RMKkPvJhLSc0V+mPyaMBg8CT
AxnOr4wmidbhMeLyByONClMwjGy3UFzy7bURQd5GBfRnj3wu12tiTGHPvJJcTDaSI7xfwwZmBnhH
Sg7T4tBb87jLnylE8UU1kuaeSyRUnQ903RW96NhoETl+2KPaGV8RPeKH6TEtlM8asBQQsiLfDwPf
4KR2JlxbKzwxwtHnGjvZE4/09PGGtt5BGwVM2xQOsEvDWdZ8fGdAg14/SH7nsBUJ9ZLn1CiV2Qh7
XscTjEtS8i+xG/luYlB3as6zG25dkVBJDE7OCki9wKLUJoP1ReKDfFs0/tFXyKEtNDmwhlwH5QOf
0l+lp50kmyPHU4a86NOpBCCFeu4LdJJtCSXEoyhYh/EiHKt7TyT295qElxlFNlWEqLdr8+OUYufN
VfUR+blowycDD7FJ2HJ9lAZ4JAjdpHBT70RiORg+pMD3DZxKzi9Eb7cFm9k2MONkZkxJ3y/ncpPo
UI85vpHsPk71WuW9zj+vaRvtfpt/xUE4Cz1kIi6hcD0MBZPguRd59cRU247WV/p3vEwhC2yWuQTp
cDAPjft06izIFlaJrE4JI5k7as9/7TMXLw2reUIdbhk4BYE0+hA78qQKO79eHVmZbS33ct2IOeRJ
6SdaZfqMbAnJah4Zh3ieyQjoPxEfsWrbJe9FZvWyRpb5ew8t4oUCpiw23/YdqQsMaJQtws1dg6EQ
wRCqeFTUrddrQiT996m/vH66cOetJ8wjeVS/fmr9YjtDKLmCegI1D5hHERGkjIobzOFb4jEBBCFp
KKBtC4yyPY0XcwevOaq1tFAZmcdPlgPTSLoc2xI2bHZE8nvhJ68Fanevf2qDaWbKi/xAvr6m9WWo
XpC0KMdQzvQVvdDOnujB/qdw7zIr/Sy/GZzmzkboNYcoEti4ga/sWUer6jtzIx0CIZuOZy2Cww4y
Se8lBwgoTvHPB+hapJR8Fs4mYVdbgdwm+PVMy1KEVe3FIfChn5UQfTC9nixaTQezAuTqhjTPQGxL
i44x31AG1rvle2fiYfw1QtjHPCLKmDp4oGrhyNTjZYhj9wZO7NSLzWtk5+ASKqlGBACDnjGs9N0B
X1QXDUaRvWBP1t0oBBpce22UX+e8DsE7ryiWuFv5EgKLvQ3/AvPsA5C/+stqQAXA0XMKZGh6hPwN
Sra6kj9nMrsu2UGHOUBJD3UOpkp5+w1sXJRnfjuXAeAQaXUgiiFnbyZQyim0yLHikMs1bdsFTBMp
6jv0zI3KcKd1lrySCAOtzla37BA67M7LQhnIGjbVpy3ltGTufomWoOlRrHUFjvwRMcLpRstf4YiD
D9l9KWXpiopUnbcnDrsFs5JRv+Ayj0CnMGc5RDbvOqTx3YPFyaGy4HC0Z8yVudksxE/j609SHC1A
ezh4RY8pIuJ6lyxDQuaGMZZDf39swVlzDipe1xzQUZpnI5SHEVwORAUMu/1P2F93n5fdcstP2ilo
KiI0VCwz8X+GtgGCoNDhnuReA26M919m+flbMWrrY/e1xfQoR9xz7Q+t1jGrFUELCsYWUX3ZyV4L
wH/QON+TXAq/c3QUO5JyTZ53zFZV1uzp+aVHK1oNEtcVu6KjoCKAqXYRURGO+tQBOplmDjhdImnv
ndg2EeyO/MlIbmktmp9LgnkcIDRivWzoZ2TO0lUGfSJPMAl1VDxUYss59AyfPBjVZ+U54fjTTeWQ
jYIN5bwUgOFf4frkirjt0ds3J98B7g8vCmfThazthKUa9NbdEBifDBwNrqFUwRe2OSKqF0MKJ0Sc
8lI2Q+Ii7En4rLlb0VyzUdqhj23CCVSAfihvzAh1JosywjJM2u3RgLuIjllg22Bysaq/OhASBAes
LqGbZURLd+oJrKo41H+EWwWFr7iSqICR5Q2hnfe/2Qc0EPIHEEYqrshQsEuKu3KxMBZTrsKsxRI8
FYAKL8+zfz/Ci9JUeEpycNUHfvSLeHnUGc5/XI0AS/nDDc05rQuWZneZsBQ6IcirMkWGiMlyUxMD
MGn1hxazCipG5CoQoQc3rrDxFlhEK/UIIfTjbc71Yn9nDZnHU068FVoP0ISNUBxb2MdT/zkNg9VJ
fW7gaJgrDY/luE/I1tccWfbtw7yIZSgO/MvyvRMuK1JGDK1h68jH+bnBB4psMNRPlrRUK45dT5l9
GTmsh4BwIaWZ1Tm1OOq6Rkl5YnYlwQcV2QlSKEr0StWG8SXWymKt7C7BJh7DtcUM9SIZhmpsjeHY
CQl8gOQ89ze2/UTI8rpWPvZRa1/EYRz8/5wiSeBkziOAjom/KeRQODZ0hsWFO5BVRe45elU8ThMl
ESOVSzws1L2ETWcXbkpM9GAZHRbwmdPajNezc3CnihJzbiFZ43PgQofGiRTU9QP+bvDUGcViziVS
V4edrrKvUCEr6mts0fdoiabUKJpIWPFjUXB9EuEXbNyLraxTfPE1KIenAzkPIjb8Hk0i0t2YS3FY
5HhUHcYzQk+9jvoyhVjJiKTeUewrSsfvVvw5+TfCLjnDW5vH9iFdJa8sQ82/Or/OGQllkgUi7nXH
/Jql3E5wrRmlWjPb+7kqT1ZSPD0PH1ZC7mNv1niVgQ3jylCLy7SuE0607VhveoSnLjU4s+QkHuOJ
HgDxqOPueEPlyEp+r1Bl960w7ENhotCnJK1dRC4cpayet1fIc/Q8ZteC/WifU69evQ9Osu57YtJF
WxQTxbJmtPyMSpuuUvJ7qHCwUN/xghhvWK31As0R+vOXz36nXo72Yitu+38geLqar7x10BmX1E7c
qx57FiLmAMZElQW9L6yixZKP7cgy0a9NgcbM3fClTea0DG+vRZEKkcdj3FfAROWel9VapWwCsCdU
ROClYCd08tJRZ9ocaoNPztWcfobHCmpn9k61Grz9cjUTi4JATAUrKZkUEIUgV5WNE3hua4m8ugP7
Yj9RtTdFvmXcsr7KpJK6SYh6rAQzV/sRL1IkFgeE+CplMStTU8t/gAzefyYSbvBn3MMU3WSEoi+/
2oJHrFPuIkOm+YxyzyJpiOGpxCsRLzNdnNghQXC10cPFALFg3tMYrXfWIMt+/ze6aSXQKPuX6Jbw
kqGgvgVd7h5GZ9VPJoHrv7mbvCPTyAAdgskxhuMMywvt8VIUfnCotGlKzfOz57QoSXgfQ+5QLqnr
Bx7cTm0O/jbu8mH6ytfWRUv9FWkxUx7j6wTMKqePCcAflnlaEzBgLBGuwbutzBvMJNIa768/wbgC
tEcBkDjAub56RL2JcYyzs2S44BljKgxXimgsl/KH+lOO6sEm1di9Xswy/SxwmQOTJJ+l2RHs/R06
fhkvm21wR37DhZOSEOOmjmQLe026djB54NAseq4WPnnHbS57FFCu8ZFif71wg12NDRrLlQX03rUh
qJ3bg5t92kVqwEEvRcCAs/kJm5mHv6rkji6xWifNBiR2g2sNRHuzM6dZnYZ56HaazngQRhgli/yd
dustJSOu6z+Q4bGtM/HqHkWlU/wa0dOUphVaduyikocoGANaIWofW0GJhK0ImOOr/h5r83o80Cdl
QM8rGgK3IzOuFNLeMimOSKh4Qs+TPov0gn1VRzaEWIh1+eT6c3kePHhrUBWOaMjaDIFiBUq7hvj8
0MjQCrzD8AdS1TSVorq/kYQN00+HThlcVdUGUhBdXeb4niaDylsn9KsBk/ETkNWsKeDVUIC8ypEN
2U/CrBqr2yJTWQH55WwRmC/6O2i0qHW/D41USFNm38D1r2HXshWH5XFyFNAkw79R9iqLNwHfFIuj
MPmV4V26mgw3Nre492BtDc+jcdbyQBSg2z7AsqVjnnU+MeIYGHsEu5NOqIoJGMA0nR3917bJcxRu
h3JjUe+ZPW0A2Mz+Z1912JnDRNUE/i1wWXYP6vgPBEfIGv6FboflOwfQUilBkkodcaRu6RudGKrR
ezvR6tbniLWrNFnT0+VltnLgqTGuz2XaAFr+9tVe/ebUdaN6zogu0E/XsJx2TA+hCrPx5ml/PtEy
fQhYIe9dVR6jE4AnlQu4NOne3vPhphG67UVJj2/XRjnfPVSvT0uC5lkOCx4U80iicKJD39FBASvm
Y0XGkx+9x1yBjbmfxRDocfWvNzId4S7CZBqqQjCtUl8SLDRmkjLEGTj4sGK1zIhwpi5d/IIeqN4C
M3dnJ+KZeNnrndnq5Nt7tk7C9NHa5/YJXZ3YViMmrnFkRx3MVVbLDe+WNSWqQw6DaW9ocW4pWnc1
Ux0vCuo6pDAIIgL3J7vyysptO2UoNGF2EbGeEulRqAgeYJQ4Mk4Gfyi8hs2AmL8PTUZ5DlGsP/M/
qQCmxhSvLzvebYbYm0wmxjeMjJNtI8xQFqQhNTn/UDxgHcRsTu7f8oHQ1QQSJOPo6Mw9A9BLfxLy
I6tECOncxs0qOPvLr9fYiPz8NtnV/VCj0RVLvnKNtvCHistUkM/SsT3qd4nW0c+/D4AnL9340ybK
VzOTygCKuek7JsoFs5kuAhpyrcGezWqEmCieS4OOqa0Xu/jIVHsvPfLhzBLe+l7KkkszhalP03vn
QKjReIuPRY8L0hO5FmJHdjOSfjtgV6G8rZaVBc0aFleaoL8hVflK4soyU4xAtGrJzvPQ3lT0BMcd
d/CPOPQr8Ho+EamEzuAjVqKsRkKhIVYENGiYrtPcJIicVHrsWJt1NlmadWfc6GgUEtJfwueA/qJr
+RwEPoT4PtJmj6SlJbCcdLGzMJ1z1lI3/CemKtOp7oY+JK9RllH4o42HClnhAFovE9yvspZ2yxhI
iJL1TN6X31rqv3DvpRornv3NeK8yOzKOzWEBgekyKmkZSeUHCmVqrIw8uGYDmdZgtkiDnyXWwzKM
3Z6zele+tkz3Sk+ptY3YUJ97i3nGPb9dERbfW23hNgSZ77XgVuNVBnSaCc4VttpSCY5rN/W2zGZs
Y87jn2PAKtZyx7fDM1s5jXffDASoQ0h2kgNe1NdB7lc+NNB7lXobcBINJzHUUIQ4DQgWIAGgm/S7
UNgRVrO2UG/ZvhLnnn/HXTtGm9Et6HtTNNQMHt4DUI1KQZt9dOQ+Eup4qwpQelkO+vzov2lt3BLb
m10sFOeiuTueRUSaJGGSRC+qtX9Y24pybvO8pXVhnYvUDOsEYcKpMLsgMt3irHq+b8XDZIdyQ5LC
IX3phTPNJewt1JB6AIVf4nGHCQdwnwyYPH8B0IskZl0Aowzs4tVUzai1W2WYEYBbOTvqmoXoiITv
7tPMS008wg4aUtQog6NNSaiqaVSmPboxTQMkQS/p2oaB/Tk+4E+4Oo25ceCzMXnU1uHZuVhC4d91
CcPYB7hBGRCOdzUoUSELnWA7iXpsgL/Ra1fGHKLH1OQLYXOKfSxzfDqqPz94C50TGQu1wJd5aeyY
MwwhW0eQYK5wyl3uPe032wNfQ/ue6jN88C5tELNGhgeR8FaKB9Kk/OxVtP+ZZ6frpGGZKZ79iSTn
eA+VH8weaWgA6T7tLplIqrfMaobTgWOXonyVd087M32in6+NDdZVuq0Ey/g8xEwqb1CV/DszlfXF
cKnDbaT4ySwozMcIRqWaKc9jxKuxi9FAIn+1fMkadd5t5O4dPNHA/wuEZlJF+qxnrnP7zBNITAap
biDQ+0pQds2M4auIfhv3igrWjW0JuoyYoymJE9N4l/fBO3/m6jVSXS9KupFT2DiZVoSbDiq1uKNZ
NVU2MYRsaJWn3VsqNJvjkEd/Q8aIqrHaNe3dN+dlMS0DFOWNCtmSkwMVG8btSWjEkRquJN1onLzv
iPRzEUaDDWGsJKnfsrmvh3+freoBM46NutA3oZWxcI1RIoE65BqRf1cOfm8FT1bCFsX5Mlb2Qwe0
uPFym2jj/bcn8Z6t9kVxj24nrof1jr3JTbYwtFJqwZyxnIhAOL8wpKqPjCpiIjluOMHIW2Aw63Hw
6fAIXJfmvLrm0IiHroXgI1asCS6OFoy/QCIcKmvdOKPHsMywqW0cTzgtcf6+wUpHHCIpPuefGC5J
98/HxBbAn3f7dpKPbLRLqfEl0mf0w5gdwX5N3IMOr5oY3RObGxx/Y6da3PKdqSy4uPVJcc54mpmR
WrO+O9+1O9ppisSdCTgTUiSmTrL9UuwHqSZThYT8UxBazoXW7Vyf+R2RkrLjiUMkPFEPe1ZI+dXe
Qb7cWo0gpMPP4441hgka7MBhc5b4RBZ3PfQbRK/2Kj68O61ka8lmza/GE3tZplwcDfcI/uQWJ1Re
DEURSMGJjrjeJhJxKFAZ+8C4w1m00FteCoWB88BwyvHWJBCkPH8BNOl11Wt9dBFVq1dsaTZt6DMy
rOn8jc+MxH23VYTNHze0muyOUeaZwmNIo8rw2GMtvrL10NTUrgg9Q/0/sG5HZrt43Ax4tFOXdjds
zolEJidUmSRuxCsOEcjf7fNrUFkNKTCkffpltW3oBC0iftIyybQFhnNXqRt+A0WSP8Ce/2h+DldS
Rh/YNW/4lSHhqvk6Zfcid8XdKIvgqaaY0O6aSPD4ZDTeiTN80HobBuY0jZVS1nUNDdB6z+msC5zG
vkbNIauTTkvkToPB+6AxHXmydIT4xsD/KeIXbItoh8fE8zCSTtUw9BzM4NP0pQ0T8HPakNfm8Kwu
POAIowpD3LG0JJvAlcK3jZVADzBMCoKHKLSvl1R0Ouhhqy4nnCRBReYcblv+aqbCCoy1DpsrzAiT
4KB6PVIn/EAsUcwKBOtQfNkQPlCoXTqvYZzAvx3Djdh+u2bCJGLsxHmj1KArPnXEUBNE9fa0jXaI
XyKKcGQy2xbjDcCngounxkFF3DvIoc4tWSUJjeYiMowAgKNqu/KfBJybMlHNg8IRldlgiO+nM9LU
hPuL/TGD4BrrL1QCPo++PF2OFpZfNhDPZlP0hLtBjL6FU6CgF5TRZc7e9lTqIdKXGzsUKjqbYcbZ
MLbDeHFWvI2tJjcItjbwXnb8KLY43ZokgL9hbm+PT6b7JC0449wKfTZTNk+HcquOEZYegmbtv3HH
pcQl1PzFMJs92D8M3OzD4bf9t58MeDUNjG4JOg8JzwD8x6itvPzqAMOaf/S/IXf5d83g4kebw2kZ
OpLizypoRL86AUa0I3dBzP6oojeGJ+cmYOZbzPzHaSK8ZwdCSgYWmbDFoyWwx11ABoKbjlCWcRgZ
V3vVIsjR252vji608EYZ/1YLmY6VXMUewxC57UbizMgK+1MuyMu7yyvdKj3f0D866kr+dktIlfcS
EMnszLguvxlfO1sCJvwMEmajKbxB5CTV3FcLkmLbutNAtVqr40YojUmmx3jCNfRNbCoThsgIZLll
4m/tyHvarJp6jqS+NL6vURrx6lLmh/pJa7KPToqM7All82zQY/Mjf2zYPaIRKujfQT+hBdZW6AHa
tuniP8IMwJ7uiJjVjMf4gF6sLIxGypcl+1kgLH/vds3aIJj0w/K+1zwJy2TERVWPPEeufnD4uzs5
PmIfDspPJm6FdZ9S0lDkSjunmGiW1jpPLMLbire6muAQ0NmUDmOcghXMvrSQAnjb4/zdkrV4VLDQ
2Eo9/PLxtcV2g10WrFJFJjZDXoSd12YCZMGp6p+OxSQAgJ0+dzivUnB2WwR3I1IyNM0A+toPEz3G
GV8ZFMk4+J5fR67j8R+7hh8B++d7X15DNxEfGWuW09/Ump0c+yczHR4tj9vvlreQWVSFTRcsvzlx
JYVNeQUMk1t2fkS/fhewU9gBn88W1Vuf/K01pmFAmyc/Qv7FU7AUINAx54Dd96XDXuraY/aJqB1s
isHwFxL7YQkn4W+pk7DzZttu25oykRyyqz7mmp3hp8E8l3iKMLiFf7nd6/wC5zrXTmd2q7VmHxWf
kWdg402i7G+DbgWVvtWrJ0Ol7m+fQr04X76AygFoRfoYs+7TeMHcCRdbim8ufMrtjgB6ZA1+r/z4
orsDIaDSzlFbZFudiLeDvIECiU5bql/iyxSaUucoer283dx3jD9mRySHwCCigAkiHGQ8jhmlyYsP
ym85EAUbKGPjgTg51nAI0Y3jaO4m6zQloDwtmkDUAAcoX4s7ulIl7FmoXYIR8/Ab2QG5JhZrUBkC
ujW9orlnHNU8n1a4pZ/cuvX7RJViAqoztPhjn/r1eMrwg6XeW2GzhjMvZc6Q7fbSa0Ass0lrzWn2
LKajmM/xzx8h3V4rj8HfZjWmHVbozhY2CrpbsCP/KtAlLpYm/zrpVjI4YaVnXe+iZsrHy59gMMj6
2JMT4fseVM7WeunopkIEwSKxb4KHpqreeEAdgbtQGG2znvhgxpxOuOkotz48mPEPOMvhLuhyI7cD
0M+FyXKKOMehWjdI57f2A0u3+NteYijGyxIRuzDwQBKkW9z0Nn0ikpFz6zbHK0BFbyjDFNPmM3E3
UaNk/OTT327rIsBYMxwHz2BGdbMZfqxAQowc0q6nE71jaLnxiMi+k4RaWVpHIvepyGFojb19KOix
cwV5SeH5eV+F0l6SZXX8BrbieTzcXFvQ/PNga+3mbJjX67G96VRiWm0+l9CAGgbG4DhEs3javT7u
jVaAQfaHAufF9rVZIyfUI2q6veGBj0QzqNmEx+D6BmZKUMTfylh59UnihdyHyEWt5/qsCiNvmw5+
phI0eoRGmmFDozeCfSITCMXAi6CsSiIc0/Wj31980yANghepfN4X9dUF36zMmeCSZ+UZ6j+aR0uI
TqzTAkGMOIJW4DpakzJFrF/2Fzvwb8bGcNULmXCG0ISfC8IB5udT8F3oodbBQ665mbo48PbTkNwt
v0oAI3urGAb6kqEiR7mLOsyhfPrI0atOLkarV5b4R0eB4xbYCqSPdF18iH4TBFXeWMXHTdZFihC9
8lHJz2K1wmqFPhF6T0TT9UAhs6aGr4MIycqWtq6XlqhkNvLFl5xTqIOpbYPMr8eFO/pBCkz5jDMr
SPtW6UCNqMvhQXDD5tGSLTWWTsHGskziOasxqodX6pYS8rBiFWdEyUY4BjwzB9EyZxWSvMGdidQW
p2ojmz2fX6UJTqb5b2qIb9C/XW6bifz4QWAou+cRxY2XKfEd+nXiXN2Fk+n0QM4DISbVHrbDGaBT
H5bmgmcLAZPrqOjk1Vqv0tT+06k6egFAhnOX3SvUz08FkrBnfk2ROnXgxuBSDgBPuaMf9F3nceUD
Uf2BeDrh51GlvgsK1snDqm7sLeYlMNdSi2dkSMpqFKy3X4Jm1TAM1paIiyXAcimfA4igLi0+m7f9
bzMY+dh/jF3i9vB/iLsOlYZFQmr8GqFddHnczl4tEuFTEmCuwSfC9RLgXqI1OkVazn7tuGVDNovb
6hc3F3OMcDp7mOjbXF12/STOq/UsYdTf4iGZOarHyn4Ha73g10i4AcwOXAicfLqNkYvJlAdmTF/E
Ia2RlvuZuU5ypC+wqwDXeds+tTSsmOyJY+YcO1cyOLAwFEziAAiMk1fDuT6zfb2ssKyEt/C8VaiP
sD6mjLuT0ZCnZgRpyTIDgXxdp5G+YShJP21LnLz1jKGAaDeqtvtY9tRUUbJbpJNyWgie1tDCtpDW
gYZNOCA6KJQbhwamN/xe16/yJBdTyaNwXFIIoGPXUi04XgVTp4m4QM3/x3at6Ga2QFwuyek5oZz/
jkb3CKTdJ/1kfBck18/8xJb10g6LJY1j4w60tTSISC4NuYXHMtJC1XMFBIqSx4JfKDJo/cHymMXo
oeF4DeRGXlTF2fdjRPYukZ79b/+IJVYMghKfB7G471slXE6bGezAMujHq/3jfeFKmCMBh9dgE+ex
tRf+T/BErPPfs/cjMVGviQAzNFOUeZWP3xv3Xz8ZubGFF5eFjQuf8wOp9DRXfkE2HUn9eGtNMja/
T83uK+wz7eP8y+yIIPuEDT6q8UwV+nUQGn4p/nGJacHpNTwk1Ktokx2voEzAnFlI6yhSB59z0Rx3
bbmyozFucjoRKBvvSTU9khRhIjkNngo1VLOfsEf8lvXu40DoZ6ZGcXDfJd4+oPKD+4kzW29xTtJj
c5w5HIaAPXP5Ufv4wqZhGlZjSgBk050sYxR6H05FOdzEHkiPE/pf3WDUGeBwTbz77ohlFOsvAoeG
uPH6zZdS+TZeU8bCBgB3UKwUA27QVpbVwArV6nSF+6mzLYzGhdgrUneGHl8TDPklmVIWOibeHJ/6
nDs0VNBFfW0L9+GHt/wvaL+DuoTqOL9Jc0pbcu8wlV2Q31chsvKUhboM6KCIyTe/aeh7R4zjiT8W
ZGXKliWy8VHFVhK2ifi/EuFMb39ZUhHnDf5E7HwSnZYJUkbmeJ89tf5Ag+JtPJ1YwxI+Rqja3E2l
epe0VhI8fj7YUHYhroIF4W/sZRrYfCnRqc+EHhitI12LHagSKn5NXWGjUDnYftbu6qaipXr4Fwjo
pZqAZ+0nJsxmDPvmuTMuq5KzwWqO20imJGn6ws1V7qNlKSNVhA+KCMTvQnIaAhKRdoW8JBNR30yR
LNcLj1nZWQm3KSlCofOGcUE0UqQP3v227jIauED7VQtVBSeh6aAWP5yju9HkNX0vJsQFK+RIyuov
ocv4AZhDbtz6a/VDlMl5liHU7QH3eBqJhpTjED9QUdYujlryDoD5eso1p/y/JFuVK2meuGWcbkJg
FTZ4X1Lk5dmt1FWtfokDsqAYJG/P/8bqQp9lyLSXMiy9c8d1jJoo9XepTbl0R9X6DpveY3K1ktNR
ECYiJrds9WfDD5UID446H3Uc8vNgudzE3beD996x2ZJfPXtay0044qg3XdfrYT5T6FDLDkFsU1Gr
KNQW/3b3FxCGmMk/+Lp3QsXY3nfA8T2QFFc/blKi7pk8toqvOCMkRjRJEvl7wLKkQk2+LBrwgAuO
s7F6i+BhKOmNbhgwT3Wmwmfn3uuReu5LjacctA1mXGR3D0D919slh7SOIClTQWlcfq7GOQcJ5TOT
N6UcS2iZqsaZZIByaGY57fLM9YcscM+j5ubvaUR1eZyhjUp+cz44GXFRIBmciBxnPvm/R4olz9Kf
df6lcnlU6RKTZCrOChw09BHQokgk6nYm+6Y1vIsiPp4k7lpi4/tsKgagfOA9t3MIy+dLR8bftsOo
3qYgoijwR7scMFcubqKDNQzyx+dnbCiFLsQzX/R57ss4RGqAgiglqgSKjODLzqyRk8X2ITlMzvgm
wwLsxJbIv/yZbCZMI6rcaFTygwNqq64Bw8HIiCqC/oUrEiGpAKNBDJQf98+pwcY9qa4e5Gw4XDgo
mYtSu4ty4YHtsYsho+kjVrR/jSsxN0huhQ+FQIX9VY7/g0+IcJXQBVX3hlM+V/KSXvn0lKnhKfBb
Az46qnDVp8veCv7ASkKIDfBBUtjEK8hnj90ZROUhQn5MoCEcWahiuoDiRsaMbxUpoFwfeQcZtCge
5mN+SiLCFVIKm4+ZSLU8/56AfKYf1G58TIbJcq66EK91Tek3u+lw8cGBRt7h95xIaK1QJlSx7yuh
MQxyhJrZfp/k6Qc9iwMfGm6I/Ht69i1+CuMRT5IwtWu30HU9iQePfMJgO5G+YgCNeOA6oVo7hPfO
OxPd/dv/gM4hXuDZJX0dckyj7XBThiwD4fL64nh6xhUGFYNzZG0GQjtfbEWrtrPE8K/nL49HJKwb
O8TOjkj9bBNo9FWNEw9CqJ1Z4peVVcbn6sk8sTiFbSzMlv1/OVMER9Zv+MIOb/ALRE8FqUb2lXyH
Azx7+rrdgxvjG6R4M770cU9dh7c1gRS5lwglqghHRz8mSUhYTXz2utQNPL0m6AHJPsIHqtVnIcup
PyGB4AT7s7csBI8j66eBPpg8Y154DvQfHAUwyfzALD0FFrxu+eklfm19CRY4b5lhivv7DDFbL/rP
fefydICsbsKmxCyLdxdFafKHQ6iJH8rdYp6F+7XKj7GWdrUpSAJ2E2/vDqPgOO8H80wWP7Rl+y12
WtMT5lBjbN+bfOAKOLcvSAPG2gOL+r80C3Z+Vxfi4WVFWgQerkMJ+f9TzeXxMyVfW2BHv9h+aO9M
LwJadAnE6oBX1My1YHV/JOBvUMpjio9l5KthTNj+gzu2BLelsd8gQwd6///BXjvcz/E/g1EeCKjR
+ZnHQtmISoksnW6yMgCq2KcOVCKGcQts99T70BL85/WiP+LsijRJU/b/KEw/0vEe592TiI8ZLzW+
cPJYtQaTEecPt8EjX659cfHfTZNbfd9E+/6pNhsI7bLMpqJfdXadj/UW6VBLVRwlw6tPxOdzNnLh
AHWGwbWQNclpHf1xStYJnhbufHdzdlFQ/co6JT8i+64KVH0+dqshcuzl3MvrgOpygLwEPgNIczKG
WL5V0JZ+hjPsmcxTELzwvFb7LvcOPUJx17QulfFqMVdvYrZcWQl8tBCNd1mq1cIVZtKfjBTc70hh
WobdYCni+OPCS4Alv0DIHMZvkOZlutMtuhls87JWxHwyDDwk4Tz/xZVRaHfyXcEbcowbqbBDPf64
xlQIUXoV1ZxSrmcuLMu+xUKZdXEn0zyK6KnQLp4nUlfSaHYJGvLGk1XWZaBmpOPte67KEo/hVtIz
bshrjQw2zo8hGlGXQEtRYWE397aOLbQdV4YddohTrynrpPr798ZhFW2ciEcoBiit2PkEHp+0ds4L
q8ryHVfV/M6RAt+3PanhCjPDgP2w9xK2ecqvyi/ZFAxx2UzvEO+Z4drGZUue8Q1DOj8dUFYRv5Qp
xQ46MzsXf3KQaTz3cO9GpBJa5+bkgKezOwzu0YmKdLKxHOuwm+Sy3HW3XwcFD0sKj2WPdKb5ie3I
M/QIYnp3YEs5gfPXsrCACbuaf2aTIt/ykcRXQHu6iQBJliLQSoa3VeMLSa3RwLCA2bsKrftF5O0X
eIR4YtlNh2atqKOpl9NMuH1ZNsz56Jky0w0AcWMmZe/WC/GSVBpfJeCz1PTdgiOonE23F9e5I3tw
SKeIHPpOpUd5iXRKVpUIblvaAW/9Wps937YvHWjB+fS0iQ4tedqpSN5dIQQTZtR7T5qF8DzgUp7q
+yImAHpF6zgyNCjpXHAmmAYM6l1ZB3gw7LcUXZnIJGt1esHeuB7dWo1UxecgWh+wbbImtNKK10vX
eDikK37FtYFM6A2FYWugRggZxXPfRV3wRhdhDkkOQlvvWzSfPakG7GeyFsnOaZ3YHzHKJTUe1VhC
fdjBInHJLMDcyrI3RZ6Fwo/kNa1OubJ/QwdFP7r66YAUm+r7zx/9wTApnKgnZtxGJRDYrHSKPDhs
3+THISV3G1ZtnISUNmJX+7efg8ZAkD3KIlniN1aAlQvUqAFscTVX45fRBCLZFnwHEr1HWJm6XEQP
BckEXYnmBZO8gwlIyFi1PQkFo6DNibjIGCNGYIz7GMLajj/z8U9W0biaPOYae6r8QzgNRGs1l4O2
QNitsj++YjpEkUj48/cRKWJhRnbS41DXgu8rwUKBYLu6K7US22Ish1Eb87m1OEYFQiWHWoGcpIL4
AmOUcAa5lQFFuaVrakRlj8Km8Mbr/NkN0rDjdGK242aLJgzHwF/OsAkQ5WaQbj/StI8lmL9QQumN
C5SibFeUxfTFO21OsqWQH1ch5TCp4KuvKFcV+jklOVKMSKclh5mi7Sjo06NDDQp7GCjNig/4s7hH
73EKQgfpj41Jces0vzGZwpj/SdjwEPloRB5XxeSkdL6AkxjxtTMGrSAas+hzCf/aqUOTswPW7Vez
s299cRpsRKc/qTPvvOHZEptk0aLrrWo0Agkly3pq7LUAxFm9nB05FTOARHYp4F9m7DDIGvlYPgWQ
KFMQ2/KNRnbKtyQ1KkONKB1yRBRi5CXiAn0x70OaAOQYbfqKrRYqHt0ENqvq8lasSLRwDLsUhiVH
kKXqHb8OK2PzRXuMRvJCAnV7Y/ljziliyCjX9CGb4t9CebLPfwRjqhfZr8OUW8eTQ6PZbJ0Ye79k
lFKqxhKMlH0RCtWTaQGfNKteWI3+F99hYEqDYY21BEgcllD0KJzuCw89muKIzToKS50kcDqjLO3R
jJhMCrxXoYFrmVSUZdvwuztUpFxeG7F1mxYHVyJif8eYZi+rgKr/u5eh24/oIe091nFor9a6HErp
o8O4Os9gZFNg7S7ppFrAUYbn2rINGmbBuIJBmFgfpVgI/Q46dG6fX5TxYD+j/aA5BcCKHge0kE9l
792q+fzkUNKeAe5vyP2D93g0cYY3VIZ6pfUciKztd7fYCpS9XcOMVtYKXFvZIf9jRkbPcussD7xK
m88yvRIPYL5GZy2E8okKGAasrGCx8PQ3Clv1ffTN9orLMK4VJ9Dyt0VvfVc7qVXpfXIQ2B2AYev5
GvmnNM0bislsTxP0U0Ys49s5TKpLWbVOgiPPIM/5A9QXsl8n7z7VDV69ioJVvaOO2oSqLIvYX7pD
dPAJRmJ7GZVSEh/A/CdZJ2NBBgPj759mSr5k3rGrMC5tgHw7TbpK/AijW7TeRaGBQbUE+0N9BLzY
3cNPOByjdL0pWJlutBGbdhxQaCNltCdBSi5GVNzQ3hIcLIUa5AL/6zSsXsQewEOpcgWpiG5sdXn8
gaZiQA9kFl2kWsQZasxEVhEpd2T/zJTBv6VNb42w9JF9YtDWiM6vfu9dpwPjmq15GMyGHpRhDQsS
JncJkKtuOyBCh/wD+TxtR8bBK3S3Jlbbba3KW9o2gZBKh0vWhvUBfTxTNIkgs8ld1SqaiCMZRcKQ
Bcy+XEwYVSNACG+fkxwSjOgTN7QKTOt+lwcTC2oXKlioZced94U6lReUGkpKksAgF20yMVZiso3a
UL+29voSL/clf3zrsvZEW5nNZv88NCETB6Qkmha4wAPTgAGvD76hkY4V5tH7ZhAfhILH5y13gA+b
TwEsEqJmKT56mBOipJYNoPpOlE5e2ON5xVmgcs5iiOIjOrUj5Juj3yTT7j82Mc+VAzFhwW4BgHzM
Bn2Xlznp09Pk+BgnIljmC5+icijGPtHy1/o5AVUAmP+hHGRNVvzUQubLdY59xuSwCQhbC8vaCz89
v/M2xDtfRwdmybMKdsoKCaGjFJi8QC39CYDLHF7nB7Am4s+zJETeEWBhuiffMRXqj2K5mPDlRFtw
fioGRhjxT+zME3HGo+gYSPcK+KyPl4Ot45pU9SwYbSK0O9Zz3GssBJnfeajPukiZUojvV3F8Puhd
2HFY6RB8YoVjpAjJYcUbuhWheMBQvFXcwRAwgKrQ1jqV4Nh2Zxfb2a6fHrDKmNhA3y8Sk1Vyp4Ae
YkYnh8/A/Ho8IKYeMQ3U/2YqJ6whEbFa+VkVvinnneToMH6ERgSPEbABoecsVY5fYG4Zj8T5EMQb
fs86QTRjNwCS6BiIODG+BwRT//L9ER/avthpl3F27hoasIlQ/VAV4IsyhBNjC+wGAexeA5slJ99j
KlLi45jr2Wt0X/c8IXV9ehmrWkrE/nxzdqoDlrEY8dkepR0ezMn9nvHzGwgOm3ToBepiDtB2VSYm
5HTvh92tT3tolD6imK2EOYFm3GgTKuIgQbc3sJS9cqwV2ZDwgAZe4yK76ER15yx92RSter8QkuE2
F7nlOoUzn/403oKg2nezVymNaV44O7CbqPk1vTso0b9H/Xx+PBDgdLmL9dJbQ001+dDWbLu6z9Gp
iGUPUKjNQ2M8bIFc2URP4jMM21VFTzil8LaRZUZq4YMjPfNFOP1HsN9ch3alVU9jjOet/uIYOIs2
jHpPFH2tsgFiAM6dO+yGaumhig4WiixCVDFHQyGL8761DC/XRyKdtFpXxNYlLI8mdAGz1rtvqoP8
vBosIAoQY3wXHmET4/+kkG8BhXD32UBWlCnsiobxxoedsF5Erkzsf9Df2gUJeGCPp1NvohX4NgnA
lj5UGYRjIpT+CPcaQSAhCu0VSUI8r5y5Urqz4G6RjXUsNiLmc9ILDPP18DzSDwZIvyaUt+kemPiG
ZH32yjbnQDAIWd4qL4tRDYLk8RNriEesOIVXQMBaC+cRYycd9FPeNmcVWRCREf7TyR1ytMp85rq/
uRMucd2pPXM0NqbyVK0Us/1rCDw+8pt/y1EFuMM1gZtdo/dH01I4R0FJetTm0hRJxlEvd26YxSz6
TTtppdy1hzepUyJdaSPApwARhLMU9OIxwT1hTqPLaq8JO2McZjPL6mMRMtEIbj/Z5XLikpY1SllH
J36zdgxCuhb2+mx3U3R89EeTTyZPQPvtRKwWU4Fg+DCLLglZPOz7u6ZERWhiGpsyQm3IyOuVwO+/
I1kArg2fCUkj7/bwYqn0f/F5Nz9FMQCaL6qmcz/XEZuksEpNPefycpx02HOnyBnrlTBE/JMUnr5N
EPN6VtNvUabf+U8JxW3aLPXUXrwiB4vvJXf2vcCqkkoPjZdoFz0dAsa+co/oo6y5j4SdwoxbsvbB
XJDfI16RC+/ONHUfmZ9jc4eq9SEkpgLgPaxOCCXdSpBgjRsnbQ4T0pPgTa54NmJyVSKY+vQTbWKb
moQ2o1VE+aLBij8bnBrRFoGup/Q4L7GAMmzF26wDlYozaYqdCeXHanV8pxEDA1s36uQyAuqnboF9
r1+yiiFVPN4KPRtYQMjUadkkmRnXXGu8LqaU8q5grZHD0tUvzBhYzVCyg/88haebSsU5tF5GohZZ
ZFONL65ye1HWER0shH3vVjEQ4rH7IoXYfctxeTKea5b+9aRfnw5MAo3idsKGUINCl3JwZfme33Pf
kAT6rdhg9pOfR0ZOEU5l2KwVoHMIqpa0mvLFb0ElglOmgr73IMsPC3yMz8qBcOK4LyGnbuo447D2
sNi3GD3xpEf+/di0vwqEswC10GGIcSI4ESCUGfkXmhlD/4ccmHf9Oe3+253Lby7BI30vU6sL9Bfq
AZHhn05A+IArjITR7FpNrDH5TJ+DiSX2GvhmvJhT3h5D/I8X89XQGBrCl/H/wKpxBsnG0OstjF/8
DoFHH8cyi8xLGb1nncwpf5z7hpgSaRbkpvgHIB5u0dPQVt5IAEZLA2mvvgbTIvcvot0f+0IDws/0
M0g7LDrBS+epuYF3KESLKOy/jEDePSAIzlBVOz9UUKXCbVO3yXLgAYQ2JGIZZsCOntrzp9d8ojzL
Pb09/agBdIu0GCX3zsy+H9q+srJNB0I3t3ElkxnNVL4KssZWCZKq3PATBgzhMHl03+broT0ypopC
DiOw9naCnwDi0yeTmkH+mkEcri8t0ex8i5ncp0uzZOqStoEiwkUbcpeGIahK9NxKVEEd2HOdjqJ+
rw4rHCJONMcHVXExhETVt86hlnJsnDTkCNuYJmjh6dELLzRgCnUnlk9PJfCmKb2dtMLXkyTKkNwy
ue9a1wMDwTPWLBnTZlJeck/Jfe/C4RXMy0X9IRwJ6lnGgTHIVFL7hbOZKdwoG7Z6VswVQxoM+uLd
CG7ZozLhGMefrjjsouEH2+FDXAVAbq/4Rwhhy6p881innAjZAk8kDSO+RQ+UqCoiLedjxIzlWamB
G3bFkySDNwpNRl5diPHuN/IcxQzDeng1c7exFNf64HiwuOMdnIJHahOkRA51xhXqasCgXIqEvVkd
Fw+zDFQ5/qXCICWCIRBim2dkPPmQ/4xNInCHTxM0gWQfteYnjpxYoKox1xmhAi32VsCPw0Z2k2p6
3RAmBt0om+XgCBpSjvmt8nnzTOZ9S7YF/cwiB6FlLDxc8PYnscYgSvQ7kqsfpKZJPi6CMyYxrUOp
BMt6Xg7dstcFQYWDQ+zCczHNVAPmg/WXobk1FiM+gYUsJGVx2b+T8KgXWIm35GFfiFADLGj8FvgF
l/tcFA0L1Lrt8FSavwIMZMjniagSfymMPVuNXZD0VKP4SWnJ0qZe38F0z7LQwEs7n80QIYA8derB
WinwuNqrFYPxf3shpfapUdjkxWWlsa4ZjrUzegLsgfffO0Cd9ufZt9DCd+SNg5ah3Tbf1jxaQmXA
RPj0j3H0SzDxbFayar2Ql90JzwEqr/hmTXN7GM9zpnqcPYaCJ6+b1FDctEOK1acFHoq/+hfPIm2L
XsNi3InKJ8CNzlB5DHiExIaETFJdVWv7vh2zFDa1UetMO7XhGuhuwKz/xukyZIaDeTHE2uiQwk2d
8tAQMMqt60l9Ecl4I3uaSvH+1I240Uis6/8rHxX+ofiay3ekQCqkQpzm+2gUwTShhcA63T/oEuBk
T0HbO2rW3GCO2Gcn6AXhpW/gmza04ZJ5uwihmYwEolba87UWP3U6d3aKVirgR46WWm9Y6xG3hXs1
MnBJFxURxaZDS2AyUgALtDIMOjGxrSKlDKSu+rJiHuuJmrNFPC+uMmoDGIGHWnyuOAsCT2MyYJro
Rt06kU6G8ePIr5G4Ynst1cke/LCSwjbrjjnyK1RHbZKAlixoWUKpdypvS54trlfb5vnxK7Dn1S6V
S3TaJ8SFQ+xXMz9smIPdNcGBfrpJJi6dFJFbIV8PHquwLW1EuKSMaBbl2e8v8NBpE9AR3mNjg+qQ
NxKIAJBMAuc6JBmPbrLvbd5/sFTqF35FbOmcfxtVdH5AcaVlIhjZGZ45UjROFvHX9HsKPppEbKEM
pTp818VLISxu42sUPFuWG70oYSACYUUwc6H5AvzS9s7YPfVGUK0SCiadZGxaMFqteOJP5nEGDn3v
bImRLhKmZJpUigIIaEFIuZyecl4q4ZEtK7MtCvmwOE3dTtR96sPuKbC6arvJS1SAbMWrNQUjjXJ1
ojAVdqyBXvu6u2h5ggW9tRIwScNbpZJlCAV41PRIIvw1BcgesUQmuWYvzrhREFZix48tNXRmixFu
Pg/Xsz3egX99KkbIQH16EcjaMsGXN5ckg8WQ6vylldWAPxEQBDG3hk9E9xBWRy+e0nYfF4y57pBj
L0cAqPuOHOi8vAG7hpG9/8vpQChGhbddT8dvK/oEudRC24YWrJcbfpUpoMFA2eZIkLPXFbwlReCA
OL7EMRcHAHXd2iLvNCVfTh/T7URW6ZA++Q2eO9CCeBNR/AC9h+9ZBOdPa6Y9EqANcsqqZUE0l4sB
yUBpbKrASakvpS+dpj5+UVAxVVHXkHjZ3wN2AAExkwt1DUPjtdtZTbPuFi53on9ryvXEGO89ZBd6
hAxkIH77GAhq0qlEcywudrKO/8Ii9Tp+eLSRgUjNxxYg9Ym+fgKjeubwUN5t0MNLaLm0X/pXEQ2a
hWyyYxq1tfo0i3XdnQ8k4NaKLEFQASGCnBNB085c2vljC2df8cVOX3X0+IGGv4L3lKlRADMZHVtk
tqig0nTeo/xQpfo+b7CVBoS5rGwY+a+H2llDfMGV7zyF8522+/kMEVsXdYqLWqm5JnUm6q8qBneY
Jlz2oLk785J4Uhxo6yEiABLg0LKrhJqL6UxgSeQrYjcInWtyeeoytHRVM3RQKt90g6AQwp0tqUnH
xlVfeGn43/01+g7SbGTM6sntWx6isBfLojzXkeWHJ3qt2Qk4rOLvPck22QATTJ8x2fwtYV0eiEBW
pKHkCWHyqla4pjR5rrznZjAFAPwAZTok4WYwgKzQE4TXsMuDLH7Pa59lCwkXokHWJr9H72utcnGq
fVhwJcafIDgGL0ynFKH7JAWdwusgoruXhQKDRQSN48iQIbRJur3vv4HAyZo//Ea+28LbzDW9q9LB
fNV7AzAhVX6OlbAgzaMWj+y1Gb8RAXML5Vp9G/0JKvPX5DynQNDtCwkLJ4ZjQnJ0VpQYUn9BnxIm
5zKfkOS6tdi9LxCdErb1UT4hgPJc/fJB/uLGxFYaFNAFRC32hma84xlP9dUSInVOnl7D+PT54QWN
n4ZccCYoarXr52YOvE0Jr1MQnCykufUs/JSo3yguCmTSOq+0PiXtTA0ZPoUF0gHeiDPBvEL94eIZ
8mu7LyHdWCccqi46FUdirxCezIQe+xB9ZwGGIT86vxs9VzSfvwZL+EkWIG+jgrayFWLiB6fHzLOZ
rVamlUbcH9YQY5AxMO17YgDr9EQEZvdTl8+zhUqeWtJ+7E7MXezngGdCjnWas6MxGyWGbVW+lUE6
HZmpDjtBa2sfgQov0qe+hKxXsd7/hYrn6c2W5nu0ZIycHcgZT5GjeTCZ58Zv4+Hbq3qQZqB4lhv+
ALGwwW+SKuFiqFoRqKweb6SH0LO/SJdHYH9el09xbzhqcoKdpV+tEI4y7VXwhkluXk8wJtS+SILx
hnNz7wc4gxMgdpvGt5sQuhEDxyKqaUDzGOYHf8R246OqLMOaJE7H09XoGgHRDvGBde3oPj7EFrp0
1OqIZ2eFxj9zWOjQdX81TgbwvEA9hhgV4iO6Xn4wt7q5aJksEGGb2/4lfYfsnsS212L7vgCW6cFC
0nKcxqnGQd6s0h369EUtgv3dLb+wpswWGR4bZQnXQcylbIg4odC2/8i9mQ09/OylRGx1Fh/2W2P0
mGYJYXY620T/QzLbPU8sNCFn589UkZjcCGoqK7kfGP7HNymA5wNM0eOV2LfKllrf7ijcjhIwv/Er
PHo7YpC6wfS1BW7qRzS5kbGh8P6jGV0viLEkYgucJrDetUtV6UCaesTykgGqLdlPMxr82QeZmAqR
csGQGvJxKjZ6aCqOdw69dcA6ZXZ24ALsjSULe88UakTQ1hHp8Dwgqcbeow9J0ts64V8yu2rlFkXk
t28Z3orz/BZezSCuz7qXZqYF3hcLqVN3VR9oTPD2WdjMeuN+OiDyZFcKCGQqSZ+dQIZsJHkWKYjS
CsDoRbZfRjPo6ha3a6qRHGxz4/2FhOeImfmANqXxiUenDchdEvrAXfaaeq2L3qFF/rGFsMkAbX4J
BOrirWGel63NTA0xuswkx5LdfMmTgZsBmiXuHnON+E3OV4sAceZc2+fAOkFi63kDSmCOMybe+Z2A
VS60kQIzUgCL7Dwb0gWL+C18BQZjDpZjK32PBxqSte6h3RtlFTMEjCHHHMALN8I3Tyf87XZ5qN+T
8JFyBI6OqqI6oSkXyFE1Luf40V6xg7Lufxxad4psnMuKE/hQ9ZKYt0jKPoUtDMhQC7kDQTmij7J0
WdFd6epBJyiD4m7YtkO00A0xgfqfLF88WAXi3InxiMnLfs0IwIVGBlxWBhA0SXokEdwZgZkjMyEa
Rdub98jAMM/L+i8LXjuULLiHotHNVpAnV/rFWCHJdObqhFpU86rd0gtx8eBbOi0r8QecK6DYcTik
xJQkcuTfNRTvjeuHmYOvJSI8+vVGc/P7pjre4but4JmywHkxzFRnRswGFu0Kkhl0EK8yBdPYWxTU
rt8LaW0X+KBhf1l+OTVfaTQABeZd1qAm7a/6rXF7L7r6Ax1XmuoOUzavAc3IPFYQFx6ZKVq5cDQ/
cjntqdXsOnC96Lqo59wz5V3NKoZRcTOua8jSmV2I4R8RIAD9FlgLe3G2AbdTfQP4NdYiGhTWKKty
MYoLwCvpTyp+tkRs52/I/wLh1sTU+xFZCKYViXSbHSfVaiCIlkAUTmsBdomQ/6XA8Ubwjpusgyvb
QC7hlT97hn0gq31JEpyRo8u8Y2y0qkj3ZnlBpg/7MCx7thVsFesc0UwvbOUQ/u1LkuPNZ76n3XmX
4ap8nYnPxHHyEF1jwqR7YBFjcci39YiUFG+2jNA7y8EyTzBXRvhJYQAGF4ThdA6gnslI33b9hvOZ
GpizcyxqU8Xla3AL9+a9XUd79k55KCA9QQaFBmml0WnaJ7dEVHCVBY0wI3HObHMrnBi3POHou2av
8y+Yz7THgXV6LO6XefWN5Wik40qY868KLo82cWdjXZpzn6D/uc0uPZ/obBc8W3fBLTSqEMLJp9LU
XMRXOSmhHq/g3/OjktpiFLKByaWKsPFk1mge2EqDM2rHQbfcoeo1gvQngYPPMVBdYXgUAUI96TR3
kE0fzANHCKMA1WP8ew/G8TWQh+JZwK+LfSHfbh1+GSw/xmpCjeK3qHRYRaS8XjgipTOEef3nSVeG
qIMRSvfjdkXjT7RYD+MZkSw6Rny7tiQ8FOYbkms8IdbojB2kcJVwdbK7n7q6dy7Z1NeScT4iDqU5
XBF4KjCltcwRRzfcIUnGgpMlN5nPVxcLqMDU/2FIRkoNrLUevddmcE115gflphdRZBMs9RZB4qwc
0kSPAUaRkgfWqBDMb4WcK8Y6Ssq1CwtjDO2ftovFlZX0b6DPBTY9FPvLwNRVmf4traBRYXYcUN2P
2JDz4NQ0IiZbSC2+sfBoIFTdOivuvxQFNVMeV4zAC5ZtoA0K0XiM6g9LNeBy4MUaSmT8EJGc1xju
wQk3lh20R0+9Xvxb4OWpbpbQQZIvyWLbe4LtMAcenm+lGTgsmuOD0h5f+KY4outSL5c1ltKNgXAR
9Z2lCVHVeiZpWoZrEEPqssHu5JL2B7C7jsyGlhOEuuXrrMFXtenGX4/Sb76R4Me5vQ82P2J4rxDi
wbGvMn/7Wh00dzo5hCAlvwnTbINxF0Q3PqoeQel8CD28jmzxV3n+cLYiBFGa/8P77BpMhsv2ke0Y
wAf5bZlaHXnjmSl1Dj13Ml6rLFzVoH1id2OLpFhdoF21SlHiTuQesBw/A6QrFgwVN0NMfXFCSDiK
uMv/aE0lrl/twNvQq0e4ni4AfUIktMi7g4zJeF26ZlHAoqFVlBtweIYyDflkbACTkhVmMjyA+BeB
YupAvHK3j04xxOoMiv2PtwNFyKRIvu0GbhOJONbSRMfzCbRVJFb8RjtkW9aa6JjwPrZ8n1QMqNsv
agYYlmpmUy+FsYd66T23OAD/OA3hq9Z2Ditl0T7r1ViUEJxU8jfwqfj8hqG8wzL96UDsGX7zbhVE
l/5r5OsUiRaV9/VviMBWrYF0RL+yqMXyOmJpJyxds6skMNAtDKvmIPGP71fNdnCvhbxfd3fFg4SL
ZrnYpYBuNQGEg3Gh3dZ5WbJYgDZmERvuTTfb5M0GxK8ZEDPmCsKcrYosTtHVQatQq4ENPubjgDfK
UnJjug/rIjXAwY5V40uvzRCQORwvkqVzULrCGCvViTX5h0DWNZR4/T5pyUOm8n0W+K5fo9T0YTnH
0AaV/6moe0bOGtzOsESwfjQd92Ubb1PtJ3fNOme3kwrRoWVjnORHjiVLcutUwBsJwP9qFzMbnzKq
3RZXxqitJVInQJDifcbg80tEhFqc59F23VeqJMEY/ZOeN38DoEVFDFXlJUTwRNZLQ7LUWRVMIyxw
RJwiFlBrsNqBwinvosUkBhD6pTTQUfi7rykCXGdPAFo14lRSnBPPWYwcXQMSDqdVcD1+kHrhWYVF
93oIwyNc5vA5JyBC9gRk6kfV+xJkQVrLNVBRIgcr0AtdZUGga983acvzb7IYmen57ZHs8Nz7Q7Xx
sM+/bk90zENwFnCXDN6Ttjnntwn4DIg0b1vuyNHUqIacAymdIOY1iDsYuoZcEb8653Eje+Cz9rVT
1FveVRuO92xNOp+exDJhM81TzQEYeXVxZAYyIk2ZS73x3Ad0FZ9R5gfCId+Q6IzDeUznK7pA0RIa
f7tgeB5oh4jv5AmNq9Cd4g3AuQmN+/K0WiSmyhjFSelbwr8kzoyLziFVPGf3WutgZlMYre0TwA/F
0c2XOuzIyn67i4BNTdVFIn4NN58acMqdgD25j3gqXeaGeDyIyH5VoX8eRqID/HUHGG6sZOJR3Vut
L4ir2uVsgutKh3P3xTgNOXMSpuUtWUE8aupDx69NWRv6HdeXuPZLcKowQByMCJULBm87GDy++OVO
oKrkCjVir80PIcNIQZ8wjbGjsYqTqgvmCCkoojAg2fnq3gAG/L/mkYvOQChp2tb9kv0r+CEIQuX/
PHkZx5ZjIwE0oEuaq+N4flpV6ngx1bhcDll9shGs2CDsDRoIERGPlyqSu3Cqk4tQJgvRsp1YA3AE
PbBjdO4W9Xfq+t2AOpeIXOtVjFQBgJT4g3LBJG9PAqGpFxt2esUSUKePPOOxn2D2dlVSWzdg2D2f
fBXhFYtVUTxtsg4THpFyyINkFNYYHqfWUrXf47stq0EYlSO3AsqDg4+g/VHRI/WhI1Y/o3vejcug
SOAfLNexPUI+YbsMDDULTJfMx636zBElwQ+FApvu0MYu1l25Uw+Vn3tTwPl/CcCIUGk8DTaQRGtz
N7gjYYy6gvFR332fBisDm47fyu+WChpz0hXM6mUhVPkya+VKx3wEbMz3VoaZrfaeA0GDej6P47q4
uuNnTGzHZ7Qim0cLphz9cDJhq8er+ukT9MaktaOb7MWO82ogLyBbBi7Gb64rbGbEmtRbIQ2RoqFU
d0K6l+bwIX2udLAxgZXp06zRW2a3GJLtMmdkg+2bEre7zRhnFno0kvoJQeRUqTQgot4iE+bmW8ya
K0mb7ad0zXUMlahJm2MwSAZw/xT7rPL+rKekukzG6AXnxN7t1+mTZZ8xjsOsXAol5rddEVg7pDft
+u/u+bw4ERSPIhXr9hDA9xPHAgEjcqBeAxh6ni3wAPpIwJXeJ1dijuEpL/e1a7jVN7Kft1z5OtbR
8J1bNAF0OhZZAW08igtbJFFxmQ1UTrW+uCDLpe6IIo5kBMzTMwuc+TF0yA47PIH98ERdsTcuM3Hn
D8HyEFIPeDMoo4tFHUCXzdtaNWYYCzPml48d+4boF+BgmPL/6561JesnM/3IvDBS7Iss1DacGBhJ
y/K18xJEkFln5HhVFBADO8ZZtXqDu5hS+gHR0GKPLtNHJJTC/2QwfAdgawjentdyR60iNph7GQAe
XfR8HZco/Hk/78tlF0H5Lt3+O2ltbWQgmy/1IVNX/qcLxe3C+ZA/lU4I1P23LMrsO8mK28Nvt/sY
xrVjplRegUVISO7EZl1en6t/rVqAXF05Eqmvnqvuk0VitjmXG5QXv1EM6mqDezdN4s1QUb1HphAq
qqiP7tYzj7iQFsFEf1d181Uu7dI4k6u4J2V10o6ikS5yCXR7c1qyHYkLN3qROpog7DDYtu4nfZAX
G5mqVjj/WWvRLoLbMm0GhmPu50ghCCgEgg9K9orDzaizNNoKKh0VQquS2pmrV34r4QDzLGJVvnOf
vhmEsv2MZV5+EdbIWwgGzCzRU0mNGb9KuKmvMh5hl0yywC4UukXnLm9otXWhqe05kIBLQu1sZJje
wbokPFwSD3leZr9KOKD35eMZLb/GrlOJw1WfJv7j8FWczNxS7lOdpKKCDY/TQqWenVoesPai26XJ
7mVq9tN+E0P3Y5XbtIq+YM3MWgzWbBOdtp9aoE6jeeUveLCaqxu6sAbcqK6KXsrLDk8INMU1QzlH
LOGze9c/p+m4jER1YXwLx7kVzfzCdK8ZT77zY6JjOLXupqwUTmNz3et+Y086Fn1C+5TnZrsdJA2E
YAdasoe/RkGzzqHdvR3lMp78RvAIJlQ+jidEC0WbwDof9qLnYBykUcBAjfVqbvLREDjBlHRCVkbf
qYu4v6ca/IRdpwYPweveGnY3V6zY2DENTGBst7Bw3kXHrdhf2yoJDagqiD2XeoY5BHHtecDF264m
2oCtbBR6U/TYvgyQNDa6YO69bPoba+PXFJ0MUQV74+sBxFpcCbZVDWnqjpb9uDs/KMm5nJhzS80D
RTp1jYv3ahiAZVv/9mqF0qQfw0vUWjSFQhToGybA0oZ2n7u044f122uYVM7Yobbo+f/jQOkTd/hF
b0ffr9lBTltyhrhi11O99f8l7gCpW5Y/wUwbg6qDdkKWSDRU40dgU5E22LzM84eLZ81bh00mMVg6
m3+bq1yE+znhfmRFP8d6Z5cQhtRd2Q3CgrewDUO6TMKiBPcX6NMe0BtyLXcn/jRHWIO453GtHVp8
malY7iiX3frEBEE9wRmO3E3AHBylCIFt3E89GaXGv+3EjOYa7R6Vd4+jIgfDj3jpYgVfRcHvhqy+
oyFCr1TCBWEd5wQqUKLf+mu2ATXCrT7Jf/BFTRF9tNtZEV2OURvNOFzFDH2rRUHTXpQG4dh6mHMU
ANNY6G0tm//VvG2CEGp3psjzbhvPm0NCaOkTFQfeBnOghHJdpgsbiY0KbEsrmFRt66LVkYGONrrl
g/qr28dA3OGTP3PMwOxJB21C70iV/Bvj2yYhRD4JGsxm4vNCkHxq9D1WpchJrBAkX17cFcUebs49
IXhNdsStUDrRD49TD7uDVM7Osz5AzRWMLBQd7qyg5Xzb2D1kvDz+z0yOkgYJk6/roIvbnPiUzzvz
6ljdhs8NniXQhnNZuAvIqSJhcTHlvmjRJUHQxL5yQC/xuN2qOzg9HPmEp6Vvl19IELQ8wNM9mnNu
ufPz0rtxUH+fEyCOx9VRzqjOjxqDU6Xg6QpQeNt2Nn6ImLviiOHP3Aa1aq4zCoP5j3EFGAs5Mwit
snVdmHKbYdBGq3J/Na68aNOdgiP673JwF2YFBSGdXE++aJV3AHx7y4Hs54RRw9QJm3fmpcOF0GVp
ObGSQSQUdB5P8X4Xu2V8fvFJ46+AlWYlMhL0DGFqzA263JPTC82ms55PU1JdJmxfbBsM+j2bdkh/
UTKfAlybdefnQaI5Jhr8T22LRCZ8SjXpL8gzc7/DzZE0Q7RB5MkHETxxqeLQ2JbfAP8QujnIK2D+
Vgyg8WwNj5/bD0aZq4hMe2Qk8xfyg6z5DyYJgL4pIzrAfFy88x6csH75C1Z4WsJJOgvJ2/Pwui2O
emUogj0SYzWSQIXNZT7LD5vA1ITbxF3ogld9PaaKF6iP2EP+d2/voU5eMf174PlhMTBUPY4vlFrt
Hh+NnTAEgV5Syuh3vzwYpiOvkDEJPkWSbcGHaKbdgrFV4SiuBH1UgxUGy/5XLHoaaBUiIwP1yx+o
MBPmEq4sVARS8lKtegkzx0bKTRxpABfej+piN79rLLrqPcFNn/jbCiCks8XH8rFBv+BoeyIFbVbS
VP0V8Bajm3Pj0Nt6/PWh8sMDilx6k49l9N2+Y90NLn4YA1ud/txRlw/g1fdww6600bxaVRTHRrxp
+1ebnFWlSwdnb5iL+mKtKYvB+cTsrVGZTkcqgo5ngK3OdM30Lmt9KiFkFAxnJ7TQ+lzDvZqnLJG2
jvmq20pKOu7Hb6FyGrSHxJhNnjq7Hd2UrYU2DUxhs5pf3Bcdxh95jAEvBInujPigg2kpoCoKR7pQ
Cs5BJOfVCkrm809a5gFX+WGnroRWC0/A5phAn6HfP4ni1p1oDkjIyu/h/JCkmoWrMJbhTMt9OXNH
+FoAVOLqfrMUGCfz7SMlQ3hwvRppbLW/PjzyZdnSQwfbpYDWURjGpOL1CJDNWZieNxib29eOn1H1
oDdOplnZEanG15zMpB4I0WKjzB1ChaVYzn+C36O5qxTmP9oH88DowOnRbX5J2/n3e6kF0SLdOvFu
7xVv3J1jzLcST3F5ZdY8A3lC1D0JnH8SBs7NNoF1dlrJGJ+Dh2Q0+blfPzR8eA4gV55m0vtOfmGA
Erd1YKi5mmteZGk3joQxGTzOcVeRWSfFTSjquDtn76xzwepMMeA8GzS1hJJS8OUGxyh/Knv4AdQU
XqFbbwEt7tBpaQjP6JPLWXM8LIlye99KWPE4HeLd5pmjVJ4LUZ92Dg+ENv2DjJm97g+NU5c7mIUK
eXAk+O3fMgl09h+CDeTfgmCkIpjODT0Bv3ivmCZA5EU8WHQtHD7HgQEdxcIATYQ/d3ZHT5Mz5tFJ
7jbKoLzn/1LixFRuKmEwclbQYKYShMlO5atk24UFxOsumME4kMhLnq4dyVNkjCK3AgaR0jIN9ohR
I8MCb4BW49lnzXyk7ha0oxmLNqEH3GK3TJPH+y2z/eP/HisMB3QFBaWp2xlV8IzlBHYAp14RYhB9
oDy9qJNvL4cLTaFzERTW+3Hv1HsAwrT/KtCf1pojdJGuT9Fjyc00RLo2XCvkt0u60h0xU+6Woxun
SNPihLKGnAOaxv84dCJ4lweodvxDjSUoCDeXMTpI/4xTQx5d4aT8/O3oC+zJ8cZwm/Wltvwcaijy
/bth7ekzVOFVbMdUXxgmF3WzCXWSEDG5Od0VsihfKNzaGYA58vkNccud+3GlYKbDXGGdEcSVkMmO
7YcehWgwucUnEzRX0iiQRQE1RKFSS3Yb5F+AW7sN87jcg6yxRKNkIFgF3bRdYaspG22egvQ2xqjZ
JHS7x9Og10zd9BHF8Tz9ZN1Jr0txzCnznUL/ETtRM0n9DOlXK2hzTgIHw4J4iNrxOlo2kG6qGQG6
ACoYVpDVRbIa+UQeyX7fb3fc7KXlo5u5z8DyPBxAH9T11lNHOKh8HdwWtkmePpciKtGm9XW+o8r7
8t3NKjpuUL9ADXVBhwAXNyJVLtlxQ5m6bm4fMeWhTtfBYDfYtR+WT8euAqBizg6NhzUjJOtxXu/s
xjoRxTSLrOZyZBlif2AT0piRJWjBMg9yxYLGqUl/ThTSvpdp5slIa3WR5sAn1+cjXIWwrzc7+9Jc
i0Dm9mr/XcVhdhAq3HaLsqtweB+NxayZBA+TggIj8w5eEzZh/vk7Z8RoLEYD5O3wqFlRKIna6JLo
+G9P9dfv0xHSCk7InIx1S29u1Mj/+uIlprBvMopcbR1CnH7xiF+5CRmi4FFaK/f0v+Upa+zP0bDX
Ah1g3wwe0ipC7KhlmjVh2P4gcG0DJiMK8M7YJlT+Ikmrk8t1mBO14RxsRFaioA4yb6bNA3XXO6Ci
SGXsUjH6q+2RRwpykleMNPMzk7dBPhr8UKNJ/dI/j67KDS99qFN5FgsCMXW7ebUV+fbJnwW/tD7t
xVX6ds27GBVD4rrMqyU6TD/5ialjn0elrKvoNQQFYi//P3GcUnh4xI8XIL2y7unBR4MZoQ63Sxwx
SXlTRu14mW4SpPe0r3vL4Y2k/zTlRQ7KH51YUQPjckolOIBWEhhrYCOTYBdJ++bz3oaittvrql/r
c7ie9Qd2FrQt8vvmNsP+TsPo1EvJ7X1iwP2b9diRW0gyNaEA7Z4BFuXsAvSytvX0v0YcU+YkWR19
DRP1PAEjU+EWGcmmcGdSbvkVT3uNCFjHytg6BWPm2+an9kx1gY8vlcvIGUhFol6fRBVTpjP906oE
VYI+sseUQuBM5GzgfNmwIXvrIuI3LERPzCKA6W4U3Tk5pLTKyUY3NWCXnwNSmzt5ueGQ6z6gdutR
L/XP0WCS3rWgmG8WoygrJmaJptVbpTmuw73gwLRMzaLDUvuyMGphulgM12B+C2qdCZie5HA01XH9
JZ96AwhgsLbnMdYR9vPbq6r820+qQDQ5498fyxzsMgFz+AzITU9TSp+ng/lArY8fPE2jw+S2VNxc
NGqZWpP7iSxro8Wwaf8SyT0RZY0rkrg3w6+CZ1hGhI9Mj5vq1q44hdU1ASxUksV8Y0usDZLTKvEt
wthBJ/s27XnwyqSwANrV4trolzUYLH99oEqHaOZtNCPiza7lkgQ0hS/Kv4Bi09jXaUHAdpQL5Nxb
FWKOeGUV8OP6Wi4SQn6tiUXlx7aOBwqJhp+ZLN9q2+FY0OIYeT0HyBVQwIa01PnJfaOhkxCSN9pz
hMpd/iaACPfGwXNdmktX8C2yIqtMR8gxxq23d7wNxv/JR6qG+zYAYpU2lD5hRWqqhLCsPuuQLrez
XP2bxcxTgeVgyi/5DEX3VR3d//qsxOgkdhugIB9uKKqp2/SByH3ul+03WM6pwGpzxUnt07au8s3z
GzYr87QYOpseXFldsFu/rtjOjx0NVflzTUMbgrSDldl0/X2G6mAMR87BP9sXSfNMdQasQG52N5zL
2g1eaiMACNu9DIlu83RzNY3oONG2DXKe0tmxIDUDJbDB4FRey/rnbj3OeRUVjvbFvk3eIhwYABPA
w/QMkxKYYSzhkWghuZ+QtQ1iakquITetMNDtcY/kUOuTYzoRQqCYSJUzYWg5MoPcUURE/uiB92hU
z5IURn/HLzvy+HBR6I1E966552pqe/cXLxj94lFnj5+bRUq+aer6QT+hu9ziv6pf7GGSZcNZNv8O
QWtoFmNeVCuV3mzAraR8hStV2VRJr2RfBYrGQu9OW6UA6rS+QMVF5ERdWHHnDlXuMRivWqe9/mND
d1NCOlEDwpHNR3MB3fDRku45kFKTceRafEJhTkVyjQLmskEBoh01IQ6ZZDSeKZAU/uv13Ndw+Yto
N47vzdnQ7a422Uo+tWOo1VOWNT8pWsRXVw9S2xk4X4M1iNm70PnJ0jHeMuUdMdBTiPuXqBtXssGR
Z4B7UGS5qY1BRSvNecWkp4IVB0imwBooq/AKD9fSzrHeiUo+mydRBY+KK/mUxrJUrQtsTJFUwR9b
QGgdKgPVm9iFhbcQd3iz5+ImXQTzdD29ZxR0K2u8C/ySby0j5yX5lZCLIGTW0Sk6TLxWq00EPWaX
P/dL5FvEm83NlnHPM3nhNU4ESViwJ9sK9ZzsbKt1R8NCNRhoTlqQfP4TADlqe8xTEjHqqE/KXGHn
xE0uq9uFh6/H3h+s6YT9LjsuKYz9dT3j95z1QOSEGGzjZvCOvo/HUAXBUiRKMrVFrnHPfixGhT9r
RD75ZpoTK9NF+whanydPlxQO5dvRNiDFhpcCiM1AWix6cZUsb6wl4K8q6WbnhBotUe229Blvo5On
vTQYRnMifePCP9qD2rVfPKR0ND04BATjaGILh/1ZYfUChYZBaj5Mj8OyZqpvH6odhRS3FwrSQAGu
XmsBQaOK7UyeV6TcA0B6IhYefXyGQyfXQ98PuXMTIwbgCM1OVqs0420K98xp5v5T4887JcvGMWrq
WF87+egTxit1GGiaR9zfYv3fhBlyYXt+df+ad6jxqvF/BJdhcSrIRLe9d2xQHcJHR/U5COJH9LFI
9S6y+t4q44JkXwJctG1dOXm0v16kANmUauVO/Qaadhq7Mx5U55iknReogo8lSlRUWyOv7AEp5bXe
62yYZ0O5Pwj41nbL0BoIcQPx4s9PdbLco03Uqd3POVdqkQClSHG/pvu+Li9dAKvylTbCnmKisSo4
UNfxoCpG0Tedi9D1KJlYUR3FL+U995mJ67+xvjNdkijuaMVVfy888F+jcvP/8Y8cwajTOXbuOXIc
L0iChb+AWTegIg17sJMrIBsJDX2rpK9tC+m9kLV9m0IkBEJ+sRu2hrgjEedjlb01iFJv6BWQ1sle
cR0uDtcdmmjanxc9U85px+VjaJAbvc3LfPQO9CjyGfvUgbkq9O0qb8OLPHoW52FQjTLNfWfbNo4S
CPorr6n7jYb02JL4PolBXHzQhL2Mp3X9bo8sEjT2ymZwTjwJ/fCli0L8cXmkdJj9wjzwIiq5tTpn
7PXnC2EtsYx9H63eYkEb6TISh8vlTS2Q8e6rmfUz5JgwwQIzjpRgP3X7vqKNK3pukq6SLxa9osNz
hNUTa7M9SwfijXfC44mkF8TVsGPf6n5s8hfhfonBpbj14Mn3RYFDzVPV5yDsSdWzcNShHs/CdBnc
2SmiM9H/gOeCteicQJCvSJskA7YRUUoWqthKPO45rPq/EyGRGz8udEIov03annrryOLYoXrFTbVu
Ajcz2SeRc8lHQJ+oz5BuJFUlQic1gj9v774RfGvY8IUMeXgf85DbZJiwiYIo18DK7o4kO6xmZ9yi
g8r8KTNomMXIjY+nP/1UR7eKbOGIDNQKl7w/Cr9YKpkL14yf6jOYxArK7QBio/U/NO3a2SizcInX
54K6cdV+HFUd+J0MULX+AJDrcefcBAOBJlWFNQacPEOYM267jAB/4nUzT2VKOlHMHxz3oVwdAHkB
GoewXcTziiliEpJfqksll4K5Knj7uPvYa2okRDL1yO0BYcEgb2Q82sgpk0Vy+uHYM4G8lL4Iv8Hv
UiTBWP6nTrZ8KpbvqNHLQl/eqwD4Z8LX/eqfA5qS7lEpBa9Z3fAYOmGGpF+llYhx2QSD/0x7brf1
gPOSrWY203BnmR0muUT4Axa05CpW55R9O0m+ivCxTYXMX7hccDVRnq0qGJ4B2zCcHjQJZ7k2J21W
k/BCpAZh5BHTOJ0BKAPT+ZWMb8Q0xQ7/MlVbSFE9ZXQKLzBB6jvdhTzWj9DwAj6NzFJ2GG4qQUNo
8C3k35MHJsjcfyLWYmjGu7nlJJwRW7v0nNxUOVCoyPmKKHIiZ9x89qQOd9Y9ExZC/dsVpxc3SUDc
l9okUt/IjxZJgIbwgR64Oz7eoMIwBucaBOJIjR7zp/+0rjl0Lk1Zy/TcGq92O5eyhy+HTeClkdBe
BZ4G8T6fa7c78sAJep1dEImFSDuAm2e7phNg6kpLJ/lLqwVv349c3xlh8MB7tMdmNa1hl4bykudu
BTeLo02HkiKEd1/eLHyc0dJJ/TBLod8Fdk83si9yXR7UwZcBaccFz981npf7gGBooQhLiLhtZD3Z
v8VmuBKcpWvPdjl6OrkhWFILzibFASIcRo59QuCuQVuSvp7nw6wlDGCqQJh3AXWjPjLzbqLnJl38
1wZEcVznX1ukQX4U2cJVEmQU77e/CMcaoI9ilDQWKzhKTU3ISlX49jSS4C+c/SVafpFY/uUyafN8
dgqdHHxm7WvKqqNMWKGsjy1KiStWns7f0Jj0Jzjy++KBJV+GcmNpZPnfVSH4+xbuGZ3e5373+PDm
/P/auFZix9AFA9Xc7W2xP4ObGePPnR6JBu3iUeRdQXU17OCQo7T32jZlLrVPHyooBJpTpZYYxBVK
9REsM8SyfcMRx0idSRDVXBr1LmwftSfgH/p4lqxLEsPkotmKT4QCO4zs8+NVUOd0UNk8YrRqq83v
xYJxHnqrdt/CG01OPjkSQ0kAiVhiKfs1MH+77OuVrOZYV+obH2nBpjDzFV0SQIRhFMvoTvO6T+D6
lscEUO7Tbc7bmAgoZkQT+/gON9o/kA4PqN0irx7JVcdaq0U2egQggZgI1M7TaAeJe8GxBjsJLGCw
u5sgAgapLDFgUZ+mQAi5j2Y9zt1WS9oYc2MEjopoOCUYST4u1Jy/zPiYvi52J711sAUuNMSQmRQZ
Of+pzgfTrWCeJ8LObBnb6/jWCKi6RIMdkwZoWypHMz14DxXG7+Vo+z2SaemKudFNnXuTdtkW2cy8
DiM3dQJCUTi1F+rbfD1qaaY8vqvZG8Ou7CAzwPfy0GUjAvV489fsa/HdVO0XwXT0zavCXhv39k4k
GPZgHj5G/rtPMXMQADjJhNmZVDJLS3KNEKBDAjS8wfF6v5TfWuPzQ+PwrJ3kV7HdlJN1SAh8kwRq
BQtcN4o40iR6KOnjxmis19QxW1EyDcsUUZwf5a9J1o6w+EvxvKJ7Y2+57r25LpbmGWyDlGHD9icF
FbAj+FJVpu+fUpJ7rWEcPH4APf1xA768StxSm871SQAVVeLStTWoLo2oHswGN8OJYqubEoIRdHwT
9Zwc21mpYz2ackyzesp5ThL4m/RvHHw0zBtjek3cEWyl+CLmUBPWscEoMoECb6NhE4S6MOJlA33a
XxGb4ldTghvxTwGyZ0h+DhB9DNu0qFjc20HohQhTrc41TDF3ZhR09Qx4KhOUgAZdgIG9R8+mqstg
5nQR9Wm159CdAry7KKG2w/rM4k+kxbEpp6UJbY/PbM2wgVG4QHNvcfQiVYGxZD4BQpAi9+OYmMqA
ekjD/ex3XxWsI7bdvWeblW5pGkFNKR6JAO5LPqGAQxAO/RjBNafpCrslEPMVMV4+1YSpF706ydx/
vc0259kGmy4FJJ/BTwVimdGCuW1s9nssU6RFi+pM1hIrXBlUwUm/NZunpjhBgKLBb1pkIkA8iVd5
tD10B9JH1a+kA/uywa1Uy8vlywRnpcb7dPuT0WzkDcA0su/YqhZuPzvrlZP35MuhYToIw/UjG6TB
3tAebClFzgvGD7k+0e1zhTEO1PcBoaF7IJopjihQslNXLKo4bKdBLzz4vkCbfYUi9fp7+gJe4MZr
W92OTTpoFzti4811hxDIXNYIxV+P88OSoCZjlnE04CH/HtvFireZKjaICBRXN8dufbR4uSuGAW3e
gCjbazDN/XiizKs43T1LTVrTfZo8v3py/8MHwlw9u01f77Ac2NQmZKdwrZquUVrvzo14e/MnDwI6
GEWYyW7GgH/7eiNBjsiZqDX/BSQnXNoLw9i4vSXb1084Em2Nm0olbpLf1dIZqBYSQWeaeZTFQACa
QakVxhRm167aafK/WfVYsojsu2rnWIhqnfFPm3Cho1wf4wtLzeXv1r2gFqUsMEA9X4xI1dMSrgvT
TJBJ21P/o00vVRdbVpuNsCLy9ieYTP0WIzxTmDH7yjwy5Y9t2JO/TnYkkn3dcD2UWDKJXNipkYm1
h1L7WN+SpmXLbKUU3GlVGdwCgtBS8hGYAeDO4Gtadeht2zxxzp7Hb6vCjbj600aGeqv4Xp6U03FV
VPFHekfI/eDgnKbOOGe1Kyy9PECxcV68znrFpwoQOkKk9cRh0dKLfGHF46Jx1LCgDhJG2N2i0pHq
XrR6BVkwugfwNc+S0WAFE3rZU8F8/D+9bo5YfB3ApIIN+6F1dBNepEii8wDU3C92oBc5T13W1dR+
G+/uiY76LzRGHGU1ItRP34nf14RmQLGD0SDmKxxTMAYGhDwaDojZEkQj1lFfT8++fVZuahortiCQ
ARYIWH7quAZvEoTA71imExUHcQRqqNGDk9CPfz+n9oE6ASug5qXp1VKYiqL6cWzDAoakCQRyqn0T
HeeiePEnGcIsB73HMfvKb5tbSgmm/ZbuvUAxhqJyUUPlSbI+LlQNncKXvBx5b4LoIDxtPEbQq9fs
1G74see0REZut6KiNzLx5lggFXdJ/YIjKYWbtpyke0W40AsuiZnHdCGJYaPsu+0cYux543Qd5wIA
tCfULeZfUjtAL9gOtHwtru21lJiGhJpSC1+/04Jzanb72JCKofr5ghyh6ZUpZ9FKMdRxirZxUOIa
42clD1xdvhtuvcTFxapdzSKKjgR8vFY5k6bvPfzpwkuSDemebElk6jRQogND7SF1MPqnKEFy5Fn8
fu2dFgPZXD8lnajI3HnRq62IimL8b78dzFp2mwKC6lqHk9gu3u7ujKuAc1f81PeJBG4wMcsRM7Gh
i1ClYc8rCj6e343ueMPLUVbQxjqLkJk8mWfdjF1Z9kp+WZx7lo7O57ZntFe5sJvzZBn6sW70vifg
oGMO8DYkCGyogGBZScec+DoumwZ/OyGVgorl5o29Dw1KPhJ248x+6kG2XrvRRI+fdXXv5w5n0LtT
gughQUFGsjtFnxnZQsrbqouIVf4pJOMqh7CiJ+frNwOUlSwRN0U0MnuubVlgnVwYS9CEY3Din3yw
ga0X80eYsThyLntuQi+2oWBDbjmvInhgYDmfrSFCkwy7gbO7lswtlrZi5guZC2INmEknwWgMKqwm
9m9evCKrNlSsNg3Q7uBKNyc95skGkIydk78LyT/xskz9d/YpM6AHOyN06wa0U4/PaypO8iXfc4Y9
kdmVLASa/23dX+NefXT0bE0o2z8voaSwzzXlLTCoGUJA9hw3dNJhu6Hq8J9eBbxAQmWPXUj/wHnr
daZkkPknH/TIHkMBs+vCle7v5QEf0dEqVcnRr4Zd4hGdye6swgy15ghZ6HKqkBPFYx6WFiIxUB7Q
rRjcibmYMZ28LXPBC5liHvyB00paz/AR+B1wLRDzPjEAGyLH+7KEurXE495wAjf5GjMyI/8oGsgi
QkU56sBAErsaNWkYCfTh/XiqOKM2Zl5O5ztgwAYf4469JyAWx32BGt5xsR/DJFFieLrhShbWqsRT
HPllY/9Vmmxo7GzhDLkSZ6UtuKhFLCqVDvOi/a3PueikxIL6T5HcKdZQetNWarOfXx/YyWVRLGsW
iT/wbSdNHqcwRMVqvzVVN9CuvzhXqKfMvvj0/VgtNURHP3z7Fiwz7XM52vU1E9744s1UB5j1UeVR
k+ltjgUx4sB8DHTNE+KgNrbVQjV1YxkOdFHatynqkDm291dzjsUqCoX8PuripG6yIHajKl9OHON2
/+57grbXmRbDjoZT8N7Rb7gNBD5KvICAeObfDI35Nuf62J6rXRwMGUxlV0SjfXxO2V+HfHgMKGLM
QiAa0DXFDmlDgp/uYoklMRSiz2QAUV29p2IQy4/P8wPFD+H72aHB88JC7TginjErG6gu61hwLNub
1X5sNxvZGYmIOyZ0w/bQ+yjJRPZGHrRct2Hh18N1vMHvYfdKrNYSV6L3WNOJD5F1y09CzJMrUWI6
gHmosOu5b2Ly5g/k65VcGbaZqnvhOuRe337IfN/zij7KnOu5y1GJEcnwUCImVc7DMUxCJ0rxGHBg
4LVs4WuG4E0L4N+RGikb6GFDR0bvW/JLQ9FkmFohqdP29TphbhQqubde2SO0V5d5fwVyq1L/MD6K
ddDX1GQq+rcV+Eu5901Xrn+euklHChSDPoFbTk3lU11VUD4YPlpMwRkgiJu4yF9JzB+xwblha5Lr
vczEJPo7DazRMQ/kxESKEzEpPHUMr3s+9WBGTlZkj0GL4ALFzUC+//XnDuxHfxTxLaoDZbbYj9Bz
W6sVBI7yxMmAHWfTkSIM1dJZwF3jMzqJUk4vBOCLdQqkuc+pkS16V3sy7u3TNgRizfPrz6EIoyox
gkm9QwSZtpdBJQcLTCTTIN+b3fNoOi8jZglyTK4ctRqsnMRw8QH+0zEd1tiTSxSsyTQBZD1PEaRq
RhquUPwoiDLZrdY7m6d2vr115FY3YSu61ZTdGfDBlAEzXrKD5WMP0+97XY8tf9HgB3/phPDbKWDH
KTq0IpEsnUVrmoADZaM1ud+p+wDGEN6nXgkRsrhp1dkU/OKzWxGu2/LeFveexKNbsDhCN3N8qDFK
66F5Mq5Nr96pYcgBAfGjh8pqbkgkhmJ4gIDNWszMSAxk2FoPcn66EdVgZytYQNYcJsRX0iZTjyLQ
XBOq235L5GOx6trEQYNiI817i5jbIkyqiafQkdDM0Wgs2el3Yg/mHYbEcS3Y1jdCNbY9148wc/7m
toDKzz7J3ubG+N3cYqaz+X5WfZYqhwUN3GxJiRsXoSK4+tfqq3inUO1m3AjAyuJkTcHSTk7aLPi1
BwilFp0fkWqBPXXm/mgwduUnfi0kThgR8GZPpzYxRgnc4MM2aB/JwDodzYtdXMbkAcCaVocdi0rR
dG2Xe/K9T0alQmhV6BgniihzQW6FtU6wuXCBhuyw9Bu6N0rZwTAVad8VbO7WQpubMTWMH8UGALx7
hhphQds5EEY8zc9PdqnpmQ3lFkwdTbLwVoMednDfy2YriFBPiIxFDB6w3Rjed5ryJtt9jR/+ukwN
Va7r+Qkm8HDZZp7rKq7buGPKQ01s8QHytfjtxwmoMez1393AlwOfBVnxNJbYhIw0D8Nuf+usJGQw
OtdTXxHfzSlkn541QuLYssb+1lbgQCREI7NvBVTAtMZnK5pepvyhpKGAG6sKVij+HieANOp7OSK/
v5BQXH6JAto6miOyO96G44VhMZyPXI6was0IFtvz42JzfBoFIf6Gz2of8BSJjq9lTj8C7fDl0ijQ
TBxD18kBroh3/vifWJyf+N+jIYIs9y7NVt4tqrv7l590SviAN7GGXRRKc4PVHycEu9AHCzMcJMut
Q6zRruulTE66A73Xm33cNIm/JfYsWeAgIkPODnD7+U8g+kGsYyh974nEokSNcyE11AZcHaIZjSGr
smtDvZdpVcsuPOx9zhnXrhkx+MFn74uer7nlIEqCh6awMAXFmOb/e3NsoUHvUMwjrZH2UiKYrFVd
44N+ofnDGmyohqlsrLnw2mzsG6nRNi3l3HrP+BadZ3zuHKN4VQO/Hzfe7Nr/+BA9sqplvvAQR1vX
Ihr8EeBBLWbhdPw6XVBIll82GYdwZlvN/6j9XQL84Df3A+w0/AiU9gRZ0Bt35xyuQy6/SiLTPgoI
v04svP60EIHZSemIab74MpHu/IbVV7v6mRc7LyBwcNTbm7A/njN3+QbFMKw62oPSWexbQh84E6z1
SrpipvmpGMWBI/6nRfuvmS5oyk9hDkoFMI86O7ilSikHMdoRetJ61hRViycJooPtVi3HjsaZ/Emi
bST+VV4cyBWNCDXCcBGKOQ9ZX5nFpA7jT3CGw9Lx+X+mRxTqQPZi25cXHBPw2lMXEiRppJrz3kUa
DdjTXBOiKInuXUqLAfiDhswyGnWD4gJi3bvEpv+FKHXRA2BiCVdcNiod5xlb0znMMjjUaf56YhXr
O2NUl0hVtYD6T540WsGFnTwPpsKRlPHrN13Zr7en/MvdjUpw7i6o3enFxEvSBbOBfx7ze8lIs0Yv
irtqmQqpcl9t9N8v3b0/NfYJHYQClLe0F+3lWJUUQTwdvkPIjrFjQv16JIdEOnT+8O3Uk6QEd5sP
ux8rVErjp+cOMSaQTSOmzbPo6E9tJGGZXxZLtJgqyG+/b6XNX2tqDTI0eNPVmmFZ4UCtRow88cnt
FW1tO+DvdujJMUraapIi0fQcH3fijPbAhU/kH40yArxOgxmBqZuRZldb/Cj0EyX3iDCozOeCHeXv
pTi21dklE48dDJRFDczl6JGitkCpsgpinhS9d5c7B5VcGM7PHEm2rySQxT57F1BUw/Ne5MLKHXLv
7vcgcbtTA/rSBgTMLQxNJU9h5iyE6IwON72BatWoqx4CDFIWxNqkb9Fxr0rcN59itdL04Cs9/xTO
rPmzhwNGdA5MucqfQddjweQUFdLZOmPB/u973cfQePjR3Q7q7mEb50Ktr5ZKr8ecEkze2cdy7yjD
3q06E3scrtUOSpE++OrtYijswS5iTbMaYgXLCSuCPQv4v+8WWsIg42It59wb3J0S3elcN/6gyhPU
hedARR1EstApMcMCmgg6+hN8ZhpOiVgZLDoXj/FRyiKe9wA/LGJvRejteeHfeFeKbSKvAq+0SD0A
Ecl4g6k1VJr0DGw5THBM2imdS5K9PeKvIhLNQ8YakBWr6L2StjoQ2ssnwL9MPmOggeS75B3kGB5l
A48dzkcdw54wNlTHxpW+XvvY07iU/Eh9qQikD0s6Unpbewp9e7SNFDpuBtKPIKiX6obqrvuyxzyY
bEdYphqpTifYTj3N5Yoa3Gx/hOazd3lSY/TT/UGM0VIUiePFYS7cQ6GclG8dS/ToBKbFoqV2rEb+
Pf9wf5Ps46bY2IQrUGOCISS/H0YhVv/WJPwvyeRLGN0pyw5oTV8YmJqXJ0dO4tO4tPhh1Bz7apEL
vvG7F9h6fC6dWCXzznB+75zVa54bZLkzZevciBSgwSSRplbPA1+nLME62tL94YO9s8M8/yZIh2+E
Em/kJORmS6iK8c/3No1ECUUA6wQRBJbSWbF717x8NFIy6P1l6fm0EFXK5Q+Ms8E3Gr+gorc24YM3
QKxDiQRNeejHdwVXk/poR8qVLrKmSeiRT1LxNu59hvKIpUo2ZtkhOKByG4bYjkwqT+rHnAlPiScW
BVgDeOfGuL7PnD2eMT9JMNILOTy9HXNx10gQnpeXjin15+89To5rYw7b9Ph/d8EeuhfCPJ+lhets
+h1NMEbNoZe+qV2MNmFAa7e+bkUzocizjClCtbmFtLFRvR56RGCEGpFoHt7/yk/4YkNuZOwo7N6t
UM6HnxMBUhWRxhxjzXO4uZ3Tptkc+pivfdenvyLjJgcsp+xmbpqKNU2Dy7CtKIVkLaGQFJnJZjHN
pBuJe1w8OLGEL2PHdj8FGeXAQGxLjXwKt4UVyI6Tge6vCQngCupPXKhVi2INNLx3gA0jhaEbfVij
DCMkbONZREn/JSxwqyuq7wazzrMQJcIjwAcWdNE/4s6m4EbF41MnB6DV9sA3kvJTcMgV2xBJvKmm
5Csk9SCZJaFkec4Itb9IsyNGyPRoxm73TLZ27eYS2N7lNZOWKVzmBDUDlBDIxZ/rWQ4P+93VM5TC
HQaIGIyO5lBqHoa5xpm8KHKZMdt+DVAsfcRKcVvfhnoLOemboI80uFsKJ5yebNro+bz4jGwcYBxw
JG+ugxCec+Gs2roDb72l07rlGky0nSM+rc1JHXBYkzJ+gvB5Ye8CPl1DyXEe8FuY7o0RLCdLS4gZ
i+f1ngfYmwhCFR+YkFmyi9SYOAzBwph5/KZlgDL+SwZwuO6PY6+fcXeg3foeWKQJLNEBoMQ24zmV
+QtWeYWE2KkdigM2djdXkc/OnOJ2fU79HgW2+3fYb+syc/3C9wS9h3bpdKjxbk2IkD663GZDIhG0
7NgYIK+Dg7BnnI3sSw+MjP0otI6xrzd/DZ/HcN5o7HyFb6MIavld+pJ4JBp/T2p+dhmy1adET81H
YHjdnbTT8LV6Jm2O1slFEPj1TYuDLOFHl3M3NgUieK6fa5/+ArzwtcGDN1eiQLExHUOd5LL7U+ap
vvradngO7CyVJnwQdlzyMxETKgbkzPPujlrszDCKLra3f3krAh0EZbo4ZUxrqGYpVzxgAyJSoQ0F
04aayui9JMhwZ7TL6oS1eOs2vs+MzGhiPfnwQXJoIi5jd/5tFkFXLHQ1GN8YVnlIxH333Wnek/8L
6dEvBREa+7Uoin+VzB90vJJif72B2zqWa1O5++G8EejF/BTZUbsXAtVKb0/m+3/k77X/knEIZ/kR
Nzqc43IpYW2eWJySrmNdZbuzRFJ7iKMAhxW91Xy+/mmDY6tZB3Kw/uHC2dBolXOGtEmol4d9BRX9
Q328HoIpClpV+2+/vOf35FSvwCbaG4YK/z00YhV8jjlX79q+tV8KaYtLY0c3t6JSKYrAy7lZ0zAr
M0VxrYFXOwB9NzSUtQZuS8TNacwoZb27n3njVFbIf1lAMCmtcH30A1JfaJ1V+Rj2GmbdNUBLB99d
JS6x0yctliqJyT9jJEqUkbGe02zobKDgbwn7TROUhforpG5x+4nxk1tJyyGepzcuwlZBc5480tq5
dof7tdDT6rgF1WDd0C9F2Cd1qUJ6nZ6j9Dh5hahwVi78dJIrBL/IBHqIzl9qRbcEd1JRC1FaqVUv
jEyF17au8sshOqIlRGdS0KwEXurg+ujbBIWv6BMiSmwmKYLYGBzcS/dcAU5kR+9YhjjeIiOHNFFM
TIcirc5glOyOWmxcSbhJYbfY6jTyV3tsI55JLs2eazwHddIbmeuxSWqzKF3fvy1Tgpz4nZbH3m2S
wPyp/+JJg7CjLmu3rFGufJqY8rUoBUcrnrnwkybhiFEt3s0iGSizrSU9Tz+5SbmUDrcvVETWTpxc
s29zM5qTJdY2DBr1w32Mkn7Y4e0PoOez3eMs+m0k331GuAepNXkUNd57dQkAjSX2RVBAgQpXZXSj
sfPIjaiW7J3k38obSRlDpCcAQJlEreG/kx1FmHAC0ffuEVq4PiCoqLyAFJlD7mnS3sq3f/76NFnB
yuVd2UucGgFjCZeCPX+nz6zqLESSPDQm36NQsAqCluw9D+J4+TLkgKOxLTh5c7Ok6JhbJK1UPZ8S
vGqX2rNKJ9H/gJfEXR9OfwwCj564yYw/QncGm+dTC6Y24ZVJWgQcOr8TYWoVdoAekGh008uU+Or8
WIVq9XGc7vtFd2ICf6fpf2X9D/ueiFt4R7zFWpcYfh1ut+vGZH0+OFq0xtZfPkVYYMcd55p1KUpd
nsGSSPaTOhghdVw6Wi4eN6j3cyF7HFM51d7S/VDi2aFJye0iFW6S5qmhpjt0wy69Uds+aGVYzaLz
xz9mFFbD280lrhaFeU2e2Zy+4DkK3+hnzy5kbcIVxvekLvq7TY+Y+n6XzOCaRrwTFlR7OetlXEC3
dJykDLWC193r+t1E6AnjzF4Q8TuBFF+Mdg2czQmuolhbYOrvMUKjnT8yIKapLtJfKc/aTTZMByVV
HnwLxZXKz9Tt7y+RNQL8FmWB3oydHhziGd+b+dmbFMobnAMlWs1HFKJPMO9Jf2uwWeyNFoErk+uR
tTACFJVCoCgObShvLCFyKoJBxxIRu+7coWI9ul4DBfj7hPF2h2XhOPbTpiK+odFoF1NAF0oxrQgl
dN6cCT7/wZ6NAomb93KOUplYonrffXt9BZCHW4yAl2ICuK/qv0F2gSKTVuzV4jcqLl2Ffm09JBq3
q7pjQAYAu7tI75AvJ0y/EATBqXAvvcI8tzU5KkCS4J2Rnaz+Je977sX1R6SA5QJtpinb/rcfuxci
cc90BtJnO8eUFICKl9QyWe5z1gyyBDNGqCFZS7vNmG18uBy1ggaOaNM3H4v7jdVNH3FqxuTtjT8P
XBNiZHg9D0iztXYQ7ldeJgLN42Tfdl6W36fEwyO6c1phvPhlJVZD1Z1aJJd9Io4mmQ61Lmrxy1E9
phnje66oIdqBMfRTKReCWcgw6EZ7Xf85C9dBIsIhlnyz8LnuQ4/CvRLZhcN6YrJqqcs2k4s2Iz6p
BWGv7nYV3gGBkPENRChdfjq2cMmhjK5zOFUjGwzt6Ljd0uC9vhnJtS6TNcSja6krtlfkHxKEbcck
gBHYbd9YSKexpvAeKkwWyciEf2pHd7N3jQXwgvYmlo/t9Odqz4Qj/PhRtjSIAaPZNIRVcXCg9+jj
nPgEYSikbQuR4dpn3iifl4PcKA7XU42F/DrdabSpwg9htMIpaP+I9rUybESXu7q07du0eBWoSKZH
oVe48tvi2M89HfpKfCtfYXxLGpqGK6ZmDhAMYzMCF9HUvrxZIi7d4UZ950jYkdHtOpuagD7k5skg
DnlIpqlk/MvRQB1BzJBoRVnoIQntxeus/hrYUUsewF1RI1jP0ky7Op2cl9tpDw7cd0zoOPBKZTSs
CkPFOCATDFB5SbQjqJ6C0SUSqExsV2kqkBQcXfczceT78ySo9G0V2zh6qBDmgwabNkvo/ew61IXj
LsXjFuoC10DaYJirod6mC1jinyvqaF3ADV7OGyiOR4wxpA3UcyfLsT75U3roPafKLGjUk/Zot+gx
Z2vh6xeBtcVWXeEnK2h26qSwBrqxyIk498KzQuau8M5e/QUsnf3eOIAOfUBybAaHc1ctVY8eXGlC
BlHVLg3s7kw/dRfzdiH93n1KQpVj4/yOX761sRWyIlbbf0UCjZaLDiREaVNBIp8LiphsyGv7MLT3
QaxcQkyYKpEEQZaPY6hQQE9PnGa6+hcYwSUfY7NQ6CQguCe0cWKavb8TXpQycr/J7vNn0bmVqQVY
poPSArxS4rrnIh7Rkx4lVsaAgBqEGAsh3Gis/mQ6wIfdUiF9eOkIXYtqw0NjxVojr09xMgbjkkba
dmTfXkdR8r3JbclS79dOOBkgYEhG7CQaNY782Zm7IvsHjezjAWJcvR+PkYh1hdqADnkeMP0Sawxa
tKifbWiU3HNpoGgn37n+ePP5HpqInu4gHHKAEopToUlcwKpPnDRi+eX0mpJQSDyD+vISJiUZxgI6
S+NDMSJ6FqiCFSeN0WbxqJYLqEG4hmsTMkcjyYKzmE8vyXb/RixvQXP5/Js97JeHD+Vi19h9Bnbn
diUxrpkZWf1EWDGeIKeBEeO0jytAsCqQmjt9kdv+eHjD9jyJn1X9zVEBmzW5yATfF0JBkdfDeHTd
/Fi0LCPlxWYqFgLxzZ/Fi9FV1yOambqrPGZK5uFEbZ2JNjPK+1kZyU+mb/zCdQr0HvUoRhQD4iPT
KU4DT1KJrAPio0oRXyxcRo6J857CHT5sRSZttY+uRWKryHMW09WsJVWVe8iPPqdv2A+r9JwTSvE8
uZU97HmPzRP+1cQQcWbeB7CdjPuKWgNnYw5B1rHGnxuRlA0A5na5Z7soI4vYG9Uf5JLUAYgfIBLE
eDgzRjSOaw7/1UsD7WReVykE0NBNsCHp8hj47JGdGaPyrZoyjrawyarkwBhveSewhYR/qY8YwRfR
AsH+3MKoQdSV6Pny1POT74NqY8M1pnSqPnc0Oq0b/u+GyTqGhTjKwVjfPJl11ofMVjPIC4EQ1w82
drWK0eqVtZJ49sUsm6MKXbFzcb6OcbK4GiSq3gCcTP+0LDcFThBIR9ngwjeODhj/U/pvZBqviHgh
ruOf1Sp+sOk9X8ccWNHR8eYxS7HnI68phbmNk1GKJGVHhq9eeGlQINUjVsTIHJcSPVXP8jEUPeQ7
sWJZ3k5gJ9xpQsYppoJkDYSuEHKdvykcWpQRAkxanCFuHhBr8OZk1VnBK8G3Fm76NYmRsuGp1lAH
DHjIwXkj6m026aHAGJs5o63V0Bv8LSWAIUD7fS8hqDMmH3QTZMNU28suxamGWKN4//7nxaQi1M4M
+7QhyIDg9L7I+m3oFWXmfXsLfjipMiWs8g3CYtcjiOet5lP6hP/tj6Mw+t1WORfS9vXGu1caSXFJ
T3EHb1lALFIT/e1uxZ13R8F8wgOYbAIVI5ELUye0t8sKymM/KyFrwBNrClZEZMjU62cT841TFQyJ
ltr409m/Fh/wcbDBPRlFPrknm0ORRO+0QveI5jwL6IP6sPRST6vF0oBpwNHPylxnxVmjNIYbxhwF
xrKpNurSCZ1L6EV0cYv7tQDWaQxE+cH/ZgxR8hgkiLZLfhGdT6BUCwjyS4LC9LFazi+d8A680zkt
5DYATxBUjsf6oG0EdBw6HYONPY3wOvhKhWZ2z5ZKWy/w1y0qofG3v3nw8RjgwSbReG1SXpMUG6VI
Mo4OpWnoFtmujVrCrfX9j6GK5pbrbXcyYtDvYUkKj25LKMa/sKm2iHj05MQIkuVk17XSTe0BzAFF
5nFJ1ImqBvJE4BnDkjHVe1mpq791DbaKZ7FC19Xm+uQQbtHvgj7osxy/XfPvBLhKKGX5ztHkadPH
hFdxR+tzUvlipse5EJ7KaUIiing/aBl+LaKrQ4S4AkEQlmP9hOBcJx+84W+btdzBkycDVo30jCgw
p1wD3i2/knaS7E3foCkYHJ7wyBkpmkjgWdjWSE7ebGI7iCEOkeokceqqusEg2kcJJDOsCnveBjtG
4y5BO9tQXoKCPHeDKpg343lcp33G8T8JnmPwBOda6bCbHE2r+834KP7JOobNlW5GZ1xY3zDZ90V6
7C2oyco0oAht0LcOrWISf/dBKv6Mzo+z7vaVMAl0rN4QO/h8YSapOi/P53bYC99ur0fzMk7VIwcG
Xdf7hBCT16w0OT4AbMJRw39N+bu3IG8KwGFiL+mLvFrrQ/sB4nE9Q539jYlUq6kyj/iJtU8vuonv
3Jn1pB+zC3dyj4HKTbLRIx3fH77fzs58SvN3d7VNS1VVYDD2qrRa1pozajN+G3j9aA2XG9Ir+O+k
NlMDC0opuqC9cDF0n3NMeuY9D9pGl24SyHMS0lqqOTgQt6USIb5oNBOao+lh369VpTis5TwPgsaJ
mQjrjZI/+S1KfUV+Xc1XIC7Fo1v8wYKhkRtOubQCnHROxFdV6M2HS7jMgganU4CKqWpSc/NkynaV
DhMALuS6oou/oqPvgDHVG2/pVVi0F7hei+oEFhaL5x9/iStJT4dHXz33v5/x50A1jmgpZIy4uMVD
E9pdpEnKfJfYfgbd+OPAgwqoxQQUudECTQWmcRb7faGtfqXuEVAwdSnTyycW/fn1L8hM70M3NbPB
q89tYfc/DrbJs40IROirEwZZoG9qgfL3BFEHRLEcO1rVWAVz7O9kM5VOZGqgr9Rn9cgimWqcCgEC
Ve+q1snZjXVuxXffmNJ7OfTVzrXgM0PFTcSCxaiZr1IFu7G9e+tVGEh1td7FaZM2TP+FRzZVzzUW
kkjim8DK3a71CwN14PA40WWPMTng4zlVYI+B743pqvu8bbaMq4TEdGlAGgHTuBjx1yoXOr63TuQr
CPDUi3cdP3y0PsRhNBXqQ6YmN1o2p+nzIVq3zMGC3mJLms2aq8gfgVsT5h7vHtmpbia4sfWUFGcq
OqkqpdueiWOlKGqBe8whYKmA5agmwXCr5HfCXcErl9nP4DJ7FgROcWh4AQcwPzn7FQPWygJ/m4Tc
Yvc4Q1ypOLNNSxTpJyqmxdBEOeFAKXapaxrFhlx1rcAQHc3E9CLBPSyc9CP6euqolus+erpz5vC3
wCq5a9AENzme/99iKiTxY45GgptRZZ9BVfbrpWeE8IS3r+VdaXtCe9lzLwTPoVvgi/ZfCM8f/xn1
ZQ23FtT8wFt3bPKlQl7Bl4J1uxwRv6IrALXB8KlsjUgqgjUPjdMmdqPMr/mG+HVxM3ZVa5aIPdel
hb9Yf5BLUXaZm7sGYChNzVQc8oKUfTUDDk7BFQN2dol4rF1CwVDMqaTXmoNXoL0cTlKuixKMbIx5
ZEnbhmcCSfyzKm9yJ3b1CcaZjoVmPRTOLyJjPX4FAccMtq//U5Xw2ILKJC57xzmQG59z1Ee+xm+S
PAlXGqo6ouii9conQLI8ao2IVJjynBOaXURfIxzU2KqbwCFQeYO07ftkQxxOz/6RUnYsaFvBza5V
mJjmDRFmDyXpSbeWs80w4k8u7jDTSBlgeenX6obKplcKcc4Z0hWoBUelfwXGGfyD6YhEW84byJRm
sj3sW4/2qoDn5NSAV8IhxhxfP4RTXlWP+wAirDuRjppL74Tbd5jPoCqDlD+1iVDtF16x0BHt0Q1S
WSRpZXrtUCkSccTovYl2WXOQ2htsnOeIBFtKwqlDlomLVB1YbxF0O+077XSAO9WZl/M2MqHglfns
HXS08r4M/jKIK1qDD69k0Dc7Yr1gGGFrgABuRO7xXHY3yIMY0CZKKP0j6Xv4bWXn1cOrtmJZJjIm
RQUlVohH23WQJ/Z51axhxDWcKoliKQbnL/Bw2nMTCBnHyD7hsWknt6cndq/MMLam8EfyDz39W8Rw
5RAMDZSDflg8jEENY3fuwA23mwIuvPxIOnRKH+yPmaaUb6p3emWOwUPeGL3MF8upfHkZ+hB91lNC
4NcmyuAtg9xOVdYfc+RTLHOQGzbM0Jt3AYs5oirNLb6YSt2+8cMXm2rlJBeuAS78+qemfEDlU+Gf
ai5dCS3lIEhUrNuDxUymrbF8TJLeCfMEHLLiPfhGPwMB7m9tHKuko3AWbwMDmI99cfJuNxYe/+3t
FDbF2r+sVEDeoJwx2trWYHXVobAfsXHTbEfvg0wNKcPtuAhziJ0EoM65C3MccwW0jdEQOEJOApvC
NdHU/nSW7UICV5mBx+rMlUOYOOj2XR2XGLHwBtydrvBqGQvLL6W8TzTjX+PIj9IlbcJWoePsIGje
DLlAoHofzVKGVVdZST1wP7Mf6FtF4eGZSWdAyV0UORWcQoHv0EQG0+pdjuGPMqqun8fhCkzrQ5DL
nVzY0JCzi9HyIt2wtMd2RmKH1u2ZNhnYbG9xlBgY6JIdVW375nvDPL2j1sk3nZW7CkjYGkxWN37R
rqFRg4ygJF5ojMljBvr5vzzhdFzTQVCM83zbcXODGybT42SAtZhupjGFTVVLW+/vTpgYKCZtFV5x
ZIY/CxRdhOWJN7ssru3x1DdYXAGFva1cWy7gcwujCsJyTB9h+IK7jvPbLoZzxUgjzeAlBOr7ssCy
ENc25+UX6WpbqCW0rZtZ4o2xL8bSah+P6tHbokxQFiLoTVYvmLya15T25lRLawfG2OoQ3z6CflmT
JqJsCQXqvCYLdDP2G1pE0ou8RoMemwjghAFoL9WjmsYhYh0soyuENSorVwAYNtqlJsSvqzggzAd1
/1knU4Nnn1ydGUXbibKRxq+NPOtt6eru0yYNPxYG/nJHIMdmhuHTFd7ktAGjQOJLGC470LxXZJ+l
QLiCtuYtZYZ3meW0Bh+jbSmOjPuohwFIl66F/8sxxoiWLArV7yVB8V/InvHb+Wb7J8KpVpB0XR9F
g9aRc4JeUF+mHr5uVBuGy/7NfP76quHJS2SZkh1SFa8wICOe4TIvgp3lhPfS7VtCZo/apaDaQ3Mk
QWj70fjb7UO44yzBOwWYKGHJ4erMGnd8MaEGi6JwFwBvD3UAGIVvbWk95tbpIEDINvQmKNaupSGc
PSTFK7cvye6zFIjbWerWccnDCAeOyCkkXi/dOplvtSO8/UeG0iFT+HTVJqHAP0cKz5xBGLqznJIQ
uOeQ+SjGQ69D5p2P7DylaTmm86XGWXeVYpPST5RgsoP2VDysjmlgmqjqHbynMIl9duR97n93gBQL
Vxjv4YwS+4zFqkr3PAlQ1SLMRmtG8+nlm1EOoPeY20FuHSymfbAtIZ/EUyzM+cDOlMZKtkmF0fa/
GNPQwCYncayeLXsdsA84xR3PQfoXioWvP8txNpaXjel5uRUzxC5u8O4RZwWb9HXBRtJcLGXmkDxp
hthShbNGiqFlGg3I26Bjb8OSlYxzXIFqCxjNajjeTi8P+XxYk0jU6aZwGrC8Kn4qOVkbu+gvCuH1
jFsEelYT2myHNCpXx0neJZlrToAhzdgnxHDqmu6EM67RJ61zv2wMEqF8B+nslgOFoySh7dvXCpHb
JQuOiysgID+y+hKIPI/utmx+joX4Mf7NDn94EWpeeu6iCEmf5Z1PBWUlKAj+IpbfOv0tn5vMcgBS
kCBl27GSSTH7d9I52w/CLNRwET5x+OzFb92YI2vTCnLSC5AxoPd+L2YJ2+sCZSlDqCedbA+6t6YX
Q1NCkDjZGbooJN4ZsR9B7C+S013SRLDmvMVpNVgp3KQgXY+DoIhO20Dfv1G/vFsl+OGwYf3x47tY
NhN6l+q9CyRCRgmRCU1SsvHExkymDRs5WVHKcVulZSK24ku74blkDMoLESrsJx+fovOckTT2ntOh
p+nCxfWwK3XanjVzjmgv2fc7EyDzCDVyV3tfQ/d43Lmd4MR6r93ZgZ+SA6S1ikeYmqXRWLlXwwD3
C4VXBce9ImN9e1cDbMLKNiOVbn9AgO6ezX1vS4QZor1CYLIblOCnly/7ZWsRG8tLjvCvQmwKSghD
nrULAAUjewH45Xh06ok7PGUgsCpXQSwLOJMUPqIw9nPfmQ91RDYfeICstrktf4UU6C4g/M0Brg2V
5lLL1ttFkHhPMpENDOoKV1L7LYl04UWA+5Gj3y01sgJfNq9n/P2O8Iea/dQof23uCtTOkHlhWMfG
NJiiPjjqPq43mXbEVzcH95LsuffRiU6c7Z5h0+UzoidlU0F5ntEmB/TSdd+bm9F1OvIEjYaKPQEL
PUSSy7oPBJ1jjSIEqktjG8Q7QohAMXbk4nvQcYovGN9pT9skEs+6FBC434kD67+me2eK+BuO25rx
vjK//Ttg9syxZ1tlSgWFYPZOPEljcZrfE/NfjPCxdYBE+PXBS3LYG3IMwHGcmkoIzi6aDXVpbSB7
V6/5JDN0+22SRs/9A3NItadVI+v6090dhEZQMcSzumVmrY93oaSs0MTlogNzWCJpfQxi8cCRxGRd
ZeCUB9Ba2dB3/ZUnut3fXxe81KMw5It9XF0QM6VmRsnML/kgYhu8UohcPDsq41CqghUik59ORtrt
vSjueSKxERwIvLStdKEPZexv1gTDVtzCFzDJ6TkgFLWmORwE1kXMER9uNYgwzY+q87dO1A2o1wgA
0sqpLr69tKVXaNRjP2ZzkNcp0uPT2ugoA3E8UrMVvxEZWYBKS+zC5+J/ccg/WiXTnkOWXJh8BPq4
MoSpSpxOFR2E83CgE49nhXf7F8ooneGdzVusnft2JFBwZ9CBi1C4wrtUxCeSS7Qjr11eDrjNFjTq
XudRbc9VWFaqoln0M3tcBdFUXlw5Ded+LVYq45SIbt4ECjmXTV2KV0JGwYrcq6hoGB+HDOlEx1ub
371KThBPc3RBUmf2CvZmF/RJw9LS6B+R2iABWFJsvlVOShes8zUUtKAbhynvG/PYEI2lO44W2roU
ISHiBCnvmqCKCjgLf0vjHgF64FGEc/idlXqgqT5h8W/9avh/Bxm0b10VjWA7NdDQTQ6DxE6CfK17
rCt8Ol0EVabOdkbxfER/RY+slbowcgCaWqlTytSUhWsbsFxwUVWAQ1v8rIejspMc4wMTa9v5wHer
18ryqhno6j/ATGBC6GZCGSzkuCBJzinP+iQUIiK5lrvDDp1BD8apzlOVngSy9+TB5IFeAA7eOUht
RWYpuHL0RPCsrdTjVHLZyPZA0mQC5nMDIXuUfPp1s+tgenx+0V3rTayBLHlK5ZZWd/9YBnhCAmjw
K97ps+4e9t0e5ukTlfVc00OcmpTxEpVZHIU0ZE9ZdThV1dB4wM9y75pCoIn0PGK/tBm7ilVm5V4C
Ev27yhKnToiEx+EGI1dM4dnW8z8P3KINU5xof9jPbWCDKEzcDRJXqBIfMhkaGamNFcTQe6Indhqb
ethIDveoqcBk+oqJSjjUijx3c0wxnKm0OJUeBEtS6ti9NXC6gYjj1C68Tuo/YuuiTEKmkWSdLeXu
x1znKvStjJgq7lOkeumqzFk8UutrhbnHmSRMXpxhYjIZVsFsoDfdUi73vquhRzniL2sGxEvyYPb7
Mb1ZPIYfvmvmVzfY8ncrw8ncSdN2RUJBBvXTOUEIOSDI8IgkbAZYhsHgKFSGKPYngFJGzxCdCLNi
ZhRUUOLUNKb8qhG5hGlQDLbFWjWQZQZfkjQqK5xMBbYxsbfZUGLA08mGlmn/OHe07Xnz7wSpsgVO
FGk7o8ICswkWKXRIQSEYqYjkUFgMzHSadvGItGnYyvPr4eVnEIh9scHeJwggqy/HbCYagXVphdko
8goF5GopUtVy4SRMwo3e4LWrwqdl+LAU41wTOIwDIGlX4SP7SpJO+MPA8nTWUTZUOQ/6O4rR4KX0
qjViBPdNFJwjLCR641kE+UZcEa79izsQjgT7PDe47naZ8vkT+eHEsJJrhb5e1L4sVZRriiu7os9X
KcxjGR+Foa5XHPHEPDtwrWMczVhOt/iw353+tXwknHchttPgYMhXZZB80q9P+uPjM1yuhWlkRHZc
YnDLYDRtBRGVGxzTF58et7mcSLfo8tJzff6Qr7KBpYm65h1MUo6KBljoX+LO+EwxY6X4CAo/siaT
tbPSxBT8YhTXHKCqAv6YGWfJPPHv5Ls4FhEI3of9vu/v4RdCQiGJUBsaEtJ9nqQV1sWKvtx95b3T
X+2bVnKiOQhiHFY/DpLCjzL8Mpm7nRwGrYy6k+oLfw0lUuYi17Kl6UjlwuS+YHkDM14vQedtWHGz
NApbXZbV+Jqy69ZhfcT876JEsmfjwqJ2Nlyai7jg35LVgihCC+6lr7mIfxkxZFMO/+sSmenzi0DM
P54uMewADIZlGafy+p9Wlw9ys1Xb1YBUvqKnKcHZzdXfoM6b86f8h4btzD5em1fFJctUAWavm0WC
axQRpgm7i72wxk/rDYaWhIcQ6yFZcX3TSxuXwIzz1Re8Et9zeDzvgaL5atYsFkV2Ll890WHYX53S
GISNnMjpDQSLegn7Oxl7JI3XTviPlLhr80I0lZFQ9eXl4PSdVlmST8STtwMva4AQYxvW+KMnvzei
PU4UarRCsUTk4mt7nHIa2FAFsBYcTY8lSOhARFkV64QDLkkrv65fNE7pAP2f4lbe97EuNYH/EK/l
04YixaJSgfRLAn9t0PqdBxIwSvnEsWgdfHkiICkVU1FnDgklKpTmtvJAL1jNgOKgdwhaQVuTzq7r
/CLnNqBfuiHIj3eHtdf1SzRsbJSGGZxWHCP/p+q12egwyP1KO/Lj1PicMBP/41L6MH0LZwCstPwR
i/mRnlkApOCRdZAPwvEIJaaITK3M9ToUIXs1ElqYn3qbv+hZC98AarF7BuHyIiIYVqecqyOiUj70
T7f4QespasewbnrQrFUuYQAe5jyr1YPweKhhs57/9StQ6XZgni+gA7Z4+9m6eZ/7ZbdhBbgYOKfO
Cnvt2sXuraqlorq4DVu4QoCk10zyW8e7y+aWATtBjS6zWS3dbbsJgu+fUBn0seevE12sWH4yg/Ev
8aopSHcUktYlcZTOeC4RLBTBL61a3fK0G/Bs4e/iC1nyAT04ZYyR8LfCzCo+fVMztycZBkDEgmF2
e3b5paEDDJWgt1LttjHkfEOhYgyTVvRpTgEA/MpwuZTAiZBG1JG/XedUq2tIJR99QWyvyEVWHqIG
f4QaKzNufMeWOvRZCbwM+pi+y5eLBapnI9OlxsNrdHvG/e/x+zwqfwbm4msAtBY10d7kfmvcnEK7
8Me32Jwjhon8gdHAG8JcHPIRuLiQa6yN9y1xhoiISf8PEQO1bLwMjlvgiK3Qum/7V0eohLPBkc/u
ShVRrgkbO2Ydbg3A37Wm9PVEm31icfC8gl8aU1DLVRESLxpGjIUmgWkzDuSayR0cv0M0RKvV5goM
iPSzOP5PrerBj+X1CGpFIl0G3143XvawgypK231yTR9Z5wvOnmPjWkyu92N5KpZwjKHS7Br55YVH
KkmZW6pTx7V6aqisoJYAS2sA68uk75/+4XXf+CmQMBA/wR9ULj5UUsDtyxK4/F9lx5cwy9irkGXe
pLGDK3ZRU+Y9ihHKmg9aNQQ6VO3p1NwypZ6V0BvEYIrbeDjJ3EU7Xm2RnL9xUseo9tA2cn0oF6C6
a2RLv6Rn/XN333aUG/NPsUVqaLnWyUg7T+02XLGHxdtHYltKX5qAEZz3VkVOSLitDvwqSRtp3XzR
yEsDN15bu/UeGzs2eoxfIpJ/pjqJ/zl4/MNSnmPv9hh/bYriLwPZPraMGD7qgkuLnWcv0UUMKE8I
UmV1NZZdAiaPNC4VwBXxFyp0IFGoGVW+xrwSCJOyEc8JqE/Ylbek49fo7Xn2CfFo62FgKfLfiaW3
pboexCzMx3dnnQHbqF09hBypyb9ryaK/qBav8hJDYtvZ1UucHllUHVk+2HxE80dVjtDMO+IW7kWq
W32UtIU2AZiAcdaEWhqx8fu5l3ivfZpBIfZdopVbsigpkEj8p1xpuk/2043ebjRSR8U55bPrgFW6
Vy2tqnhSlsJyB0odAWI9xHVHG0j9VklQG+NOJgGBKdZgo74q5s0g1+FE/drW82YI35xCyA8K8O5I
c2yodij/6472UjalTkwX95HG4WH3zsZ67M2dwwMykbMiCG7VnP2TO+f2x+HnMILYfYZ3/+IGSwhO
Z7rnnXBTCNVaUVqVj1Ej4a/K8QLj4PLlXTCTnblvIdjhywm7ypYGDwWaKB9ING4ZXaqkMOm8tCJs
jy8oLfVRNRPra4z0BTIxj0BnT4X3fQU1kbXw2PRWrx6QZLHobRjpkWbVlChZIwZqCB4guul/l5jp
NGMFItmRBjHNHbtYcnLHJrlNfnDbqEgGfCsaSQYtulwJSTQgsMcyAp3JxtT7QpJ0eJTTiKrQQ/e6
cncRua7N3KuqvjQ7JlhrAaqt+gPsMhgTix1jgtMWcAX9WCRy9uv2s2OVmNmrYpIkc7CjkpRdsoRp
4l9nJpYQddLLhNzomX1UpF6T1Ui5G3mtRvP1+dw5IfELzcs6ScOTbJFIRb3MRQyTfKrHN6p9pXND
Sf4g95MeRxQwwaLAwHZ7UfBMN+pVxg144UvOMW9Q6BObi/NMOCVpHYJAP6pxQdYzk59FQJbelJwm
lifBSksq6FsnIZYw/nKMhyyt1qpHIsIwm1XdDexYWCHxG5Nk8RP0VN0r9oWLHgyLmCBnkk6uvBDT
8QRuQ4OHD2sLW/nSp+63fnXtxmWlFF+GVHy5XXobuq2smZECBGjAgi/kl+m0Fka5wUtGu3IU1XzA
z+P+5Q/G7VkVqZp3njKYgjQFaRCnrP4sRRxOSvh7nZRcgXWhxt4JMEzMQ0n+qXNTG2KcFG2tEw5a
nVgfLCgRG/DW3DedHm8mgTzqLNkVV0xW3CXRYmFLQW0LeyyPsivw58o2YoMS1vPLcn9KSsgHfHrb
hVZ7S9osrj47OXg3/OEPTNsZ6Kfk1ZPmCEoZCtGgXjXMf1F2qvkE2fsogerKjcRDlxakVniLNS5J
monSGMhpnnwYMKCi4Mh2aWk3hTRh+kAZdQh4Hz+ppTYeesBAZKf6XiqPIDQulWiVJlfnl672n6E+
iywP5a8VIe8EtMB9o8MoH+A7L2OBnT5iPCe+MGCSe2s37oaTjviAUYzfLizLN2qY2p5MZUaiCI6L
isJ/56bd+BYuylP21Hh2U62ZxZHgmpKlC2F2gmlZr7tEkkrWt1f3TlRiWWwg8Wh66XuQH3SEWvdq
cPqJ4h+oO2KHGYKn72vz3qe/iFgUoAwCnp3dORTwH1ZKQjyec046rHglU0KUUNIhEfMZdZtvFBLo
xnko2neFQowOij/7JWvfQHewKzheyMnA2ynDmsOsOu7BVvTavUayjBjYYBR/6J8kzNsSsjwxiEJt
+tGW5bMrtGRzE3jq9kJn9SfAFv7XO0FOEUAN6nTmKImwJ9KZFG5/Brg+HkU4225JQ/iIGdAjei9A
qsuUm0EEM75j7vIU5BpA8R7eIYL/5qQYXuYLxCSTZNy3kPa/pCgpVQVTEM7/GTZZAJ9iT5UwlY/t
Ao9foFXqncPab1PI56brHRw9Zkwraycl92DvUsl9JkpDOj/T2VaLE127TqiQw3azqxBCFNfxUce0
IPOK1d72Lm8hCWrZqo4AAQLmnmL+CodVSa9A7jj+7v9KN7J78k5yleo6gKLYyp+QaPbh8/DaCt3z
z6NvM1FiB3iEaDWokU3QS3yv/BeKXPk1klMq73R4bLre92j70Q7GNNI2TG4zLwrxUt3DaOp/6GE+
sOlc6R8SsfJCrrXPO4cY9gpM/5xYf/l/eyuTho77blHZjx7L74Sq5L5CJIayObd75BausNq7eed1
t+elcku1HgvuubPX+tNkvy9/rz6uF9anEHHIDHJxkkU+klQuvebPVLdO2cMwXWL/fr5b8XGyjPp3
kHX93vKvBL+YYZBQCoJUTNrnFCKe8AgDIjuYLMlfCi2NFLrhyll6r3S5nfeep+gRGVMGa1eLNeGA
58Gz0mjoBoXc3oSdcF71uSTNxTiMjQfZTbBHxTfYfS3OteXq0sNUE2He9ZQ+5OyK0lrF5nv56FTs
90NnlCiDHBroH3cQfSm2KX2hRoXgZwXNhMmos6sMMtvx8mSv4J30/tHppI/gMNIpwOyGChGHU+S3
jqvwDdGWGFpJAvjsnQBUdC/xpqHkYtaydRzVbWaFp8J39RbqKJOF2kUf4MiC9SH74FxmGsKNk5QV
aWHCp4ZhYcOCI31u8Tm06DHgDYsT+9vBOFhQ1LEnEOdelZf5cbZ+b7S6Vmg3yWGHfvDSPj+7l8xr
wC7hW7lnVBLJaqfrJyTd2RH3vxnhRAlOhHedsXYJwTJAU2+YBmH+pAN8fVWs/ht07OFPjBTRxS7R
BYGTEIXKhXMicNSXOOjElLUc+WbXV0e9J3C0MI/0RjNm0i7ESR8XIE7Pxo3qhFWSCRj698eQk6HF
yu/140L1mRnwWNT8PuAxY2lInGGtvQqD82OPbbgbzTlS96k+5h4sKh5RgFNXstVCOUCNsHmAjnRV
MC/GO3HWPk09I0tJZQmAVxeIZBVTz09tYRqIfcZbcG9m4UWMvILjE3LqkoijAOqdqt8q6+J1CQdY
x98ntW9oRDwB6Jv+gN9GA39TAAgJgFa0bK9pW2qcF/rRGUCbgOE2VN27wYz/hXQ1lpaGA8kfnBku
MiryMA9mNp8HEoo/Mx+MeR2eMxSB5H5gkToiTXdrXGgSib0yGs/b0P2dHZ++8mH2l7sJ5OxAEfo4
/4nVIc74h7W3z+mTmApvr5pbVQXs/VwomP7Kdox7aQvIu6zso91IpmYqS6evpc4q+JCuwiqPdROE
EGZeD6PGAGIQVfATFQkob5eijIUvR9fUDPq+/kPa9Pwcbwui2FusUe+dXGkpr6mFmk2RNJIv42Rr
MW0XvOIhB35vqAC2x927PyrALE7gl7DYZp0pRF7xG0AklfwsljHN2kFMn0DuDfIm/B2mb2BtQ3yy
XAwUOBOHF46NaDeltCvJQpuAfQMYDabltX9/Bb9qhPU04ey89ONOnaC6rZcNDZ+rWb+DKHMKII8s
146DGNMEX3SHqShKRJsYGBVDE5m+mCJrhBFF/gJh8vMAPBGoju31iZu+/aQXqzb8mS98yxcz/gmW
g4H/um8rLjtC5q+pd3HPjlEZCoOJUA16AWWL25vFi41XJ33RdlReV09Ae2xYz6a28SuuMwsx5P0k
zYPhKcvRicso1Ib7VleJ+fjJrXu8Nzk7rw2doKoTJXbbscwKODZpucQEJvxZBb2apu6v/WXGc3wL
0l1BGnwwuAlj8bDnGkGL9f6g6u8Q1Adxx4v8tLBnjFwU5LB31BQDpzus+yvzK7cFQ9An3RtYwUHM
3WTQex+VQkyJu4AHQqFqI/zwh3ZcEHT2ihYt3oK5u1lcREvq77pISZZ9sijyehQ5GT86GvWLWgmB
6cb0A0CWyg56hyYL0flapKirsTVnsOcWfZafm+CBZCRs5bnLlp3bnNCjjIWv/I+pRS8KRkQk6yos
cU4rKXz+Zn6gFOMnhhHboFoSXHHZwOnDwoN9v+xT/HuxOKUPP1zVCF2y+ypQbHQinY4fMMZCmmdo
6LhQFMfBq6C+BDtFHa/rhpcihWH/vavgiLFv35Koo9ktdf3xxRX9dnq/QCnLtGoaI0BkOXLZHqn4
29j1F38PnLJHs9vcxvHbkfsaXK+ennht+uV2l7/5iJN2P9vTtJpigXPVDGHLldvrWby55oGQVP3E
M4NoG/ZUILdBzogWoekmOkzLRbb/riscZJbo99nrVazpaTfyWfW0ojuwwldVdSP5OF0urWyGE5Yq
G2SepntdPhMnaEsWr1uk/aMPMrMZ5dPoBkTG8j1eBOxAVbIHpjww9xy6mJpdp1tYBd9Kvcew56jc
YiBXAEB5MeEewqg9mkc8bGmJBVRpdhtsV3YHZYWQT8GDZX2BWyemiJbNvNnpjVGjKsCm2IdZcPyu
GHwaLKvj2+dXAMIb91XiUTLX2YNKa/lj0m0UwYKtW6TVC9/3yWzYFsJ2EUAiVd+2oPt1abJ/8Q8i
WItg8XKOUlHy7VVMx4rr58XLwOm9V6p/6ySVCmy2mw41dZ3GfTzhuyRyV5f0B1w8vRDToFlDsSYX
Cg7Dzi0IMkiRkX0WJPqmGHaEybJkx8KpCsb6BBmbf7rl7SjA6ffNim8jRdTa7tq22RD1+gSSN82T
LGW8dm3gtH7BgGMpe9s0Z/5OdHY6vpL5uiHOPjTHC0FoYtdCMwdTkFqmRvfumOtTF0vvbqpEy1n2
m1+a3W1qY/cbETMTReszAfPG6p5312rvDs3mWhXZdDvDeuWxNbYcS0gNho/+IsxXNhvA0yA3jtfP
PYUrC5PTRaZr8V6Tolb1PCYlHgGT4JWVPzwrybl8eYL2VG9/cgONvcdc8AsyxYT80dBpgw+3Tgai
bd23vAXXNxc8Cc0Iywwvmh2LJQv/Z86VbFDuY5LdY1yhEUDwdzerINrugn08A/xQBoPhjdJ/SA7j
SSMtW8tktuPR0RCpMcWbEbz/gHcHQwZY/qnJTrpzbgoalblHjOBfU4xRnIxqocJUq87f8cA3iyZf
RhMECt2x0EMzcpWdPyXtohKtIuW+E+NSX7fyKVN+BDo67n7jldLeHDXZRxCgeMv9nQRWAah+0W/B
yXg712Ld1x1viqLPOvHH6q1CBhloRRkBs2aqpXmG3YlGbSH7IY3FsVzDSK+J08MRMus6Frhf4Pdq
Bm8cQvBFnWtqsgGQsLqHIbne6aVV0rM1k9T728Hk7XGsPRiOQ2eeByfQnTpqozYHKMXFT6ohmwu4
+fznIEpMuINHOpMg1gi1IIT/AXx/DoQ51BzNF+nAQCs6i8y4rlk0rZiKv64SKtEmss7Y8qzbd4lz
P0pfziUOpiZbRUaEofUP8Oy4H8WH2SsBpajFBFE85yRf19PuVwyrqHs6EwIVCZtWOvldGv104JJD
xYtuYO0IitG1OMQBo43z01NVA/hO0ZnruyjHX+r0qpUkSaIEIhaENWlgY2VbS1Fkf3oVpN1Wpaad
uqBMjqWEPXHcu9oHjng2d0rV3I4FliF+0A97gA9T4LqX4K8synP0nzlIznOBsqy3L1+RjJHekhQG
M6Nz0WReXdGNyL6xiCFKH0iD7pKfNIhp1SI9BAWFjxIWZGoaw9iJ/8mQHy2pdRl1iRXUrL8Q9vXc
izvZP5+pmxJl7WK8oPtIwk0naXuhuUEGx5XwnJUfcVzhiPoNsOYxGGCI3YXpbB9EfDRLeHi7g/Zl
X2b8l/ntZgaONdPTkt7Juoo2m5exYPNEJ4X6lC5RQx7Y7G9Cqf8JEY8JLrj+rZ0/iiqyw5H0LNFF
Okn26lg+N0rE2Ac6gEZG6Bswyx4iPLMZy9oxQLUXXuCVSkiHCOityydm/9jRnMObPHJ0kqLDdhVT
aaQBQtQa//AfK64dlh52TvRIbt7iAsRQ3trTyXf0ZIshQnY50zPDD44YMxy43gZTqe2U+EaP01SH
Njv4XrMShER+mjbgRfd3OOyspTO3nkt9JDmWDEQvYDAUMFUTWDu+U/28LgM+v/faoHb5VBQvrMxy
SJaNO46sycNqS8Cv/zcwvaCvTh0BquW1//M78Gf2EFhgjxStAi3lUGMO9ksuP+PmGyMWoZCe2aIZ
D0NE06uihcBzgvhlja7GJ2CTFY7WzW7mLdVq3odsCuRaOJQpVOZ1aiuqthe9e5Cg0cLtZ+ulJEdS
PDiK3+3/pbOtLL5bkjj+ldAxPzzZUIZPYGmZBZHijgK1OuUuoW+fJOyv56ir3nm/t6gamfP0ByEA
UtXmD85yG77jTKKSiO/+KWw4cT3qpW1wGj5ZTOfh/NklQG2kUZN7Wi6wUq1c8YhmVc3cAix4ub4i
eHlvL99UKIKFWfNNmGXeFajdR8ZVioefcE19/tb7/h5nkCiTfyjj20pMJ8ugosUsGqikkkiCIdQY
8PVD1NBJugiceVborinyQGubXdvqfAo1OTR26MW68D2BmCoXharqOhTEM8adGqcjLPvcWRXC+RTS
YS37VGgNsVW17Z/zVoLobtUILWOGW2THEqM2igX0wINwE+dPq2OJLzDGGsCPy5V3n0GnZWplePbs
qbdLKd7hj/9PeGcnvKhTHZH7YBmhQPG08+21q553tJuRDS6vSKpAOWS96wbqza6UxQxIdPZ0UmFF
xGYLuBagTWc2OAeXdK8NC5igzhq9CYpOVPkbbNp84l81I3jEdVshuZO+fM1839dA/nWiEe/4PC7q
/ipQZ2eBIaaZ7L9t2C31pni6q69N0caUKDP7TJwvGJu9XQucbIjVBxX22tXq6c/xozyt6/MmYolO
f1mfMzt3sIXYh+a8CEx0u276lkaN1/Ytzt1A1VIivrYWq/SRuDUMhk6F+OiScUGbKPMd4Sjdxc/8
N+G4BWEe88xYzbKa2qe7pR6su5bXj2aBhpy1jFxj5rYPd2G2IDB98vRgDsFVHprzBy15EJLrnuhe
MkDDHhm+xxUK2fR90gaTfj+8e2oKmiWovOm2LBIK0TWkgCJ0zN21YKGdJcz/tMeqpXJU9tff6Eut
fTuc977lUvItpWzbCj+Gk/19CW41kHNAm69u4XYHJibO5LduVTYNX+3aztgtOgVp80nqLywRZ6fl
0ykU0wI9+nXb9jowfRCrCcGrrhb8r6sxXCOu4Zg8yhPTMZOb/EnXyhBwjrGbZGEbJsZBtvRaunVr
JULt0ZgX6catRuWJg73w+pdqhQYxmUe9NR6Qh+3BpOJI3BvwsWFzKJPCkLUiE2LBD6GVrJy8N7Mg
psJi7+Pg9dvzewDNn1LThG9M0DN004LqFO2j0bKvveFkWgK+s86xWvwt2MsrMwacCt4Hx5ugaxwf
vKVQByoQ3poRxoHuGj/nHvlWwQmHB/hcVPkJBLRGxNoh8VNJxweuBFNPFBvy4L3FbUcQ4kFbaKsh
v/Y32DYgZSGHkSt/AxJOBE0uBFsIMdyJQo1XYMX4hpQlLBWq12FSsxnQ6I0VBUOv3EnP56Q132SN
+H+O8H+P4eQCDEgmZ8tmyUet6zWGkpNfgHlJL6YU0Jcszn9i4cgE2Tqje6Y9LwlO639510u5fomS
lCP5Z7ePOCqs4zyuXF9e7LAdzyPXYKjhqedIMi6cXgwKdnJ4DTazLFOSo/ba0QuDxdOzTmJhfd6I
jhic4KzzLhDNdMEZd/SJRgVU7VeWILv9lrIVw318GQsGc+Y+J8n7ejPHXekdxGO4vX86QvregE20
Y6VPfB0h86hspzrqOxfdPywlh5cqJmub11YDkVBUTMKE3iga0FwHzlGhHSNZELr5xObp7a9YLD2H
kv7ASxiAOnaDGhNgduEnEBLylX/OQuNJGknzahT9c5o9ZY54IzX5igbxLxR3b8OQGrbiJcdw53Kq
Y3HN20buhm6QrutwMAZ4T8qlezS725F+xdouSsqWOT3WnH6oDEdKsp4aJ+rF2g353CUp1jg4pD/u
bR+nE94b3vYV3xUPDWV+erA/L3QfairNoVxoVwnKs5GdTiP9eBMNJ0wwfpU/vKcLDCy3VMtpdc0x
5fHNouaQYFAN1OwxOJE3RI6ga3OUraHeBh8sQ7/lK/6u9KMJqlKdoewNTkkL2pDGX7EGNRPZYMYV
y73u0+6UuYwzn+hyEmIepwVSqbXXRT00qfjIgAJKpTArGOcbHupwMY/7JUnwHGSlXaAeF8juV1Fr
IvrenTtlFGJrSv+8Mrgys5GBXAZdoQxOGszkUpvWctggrw2BXTzoLEfKugAvYDvgwdph2G0x+CSC
RG3cRSHTiGKKu1UydAZhgtlSroSNAeexJ0w8UAdY0QRXiNj+M66wfQ1PfEDfKCFPuvB18tKypUAQ
M2GyE6kpo/Zjig4HHLuwoKSqxlzPLEhZ+4lozLuZ0dc//Nq+c/5RFQ0kIBDmjNxyglRd/DzwPrBS
c3I7EkAp8Evu4bSJo7w1QQu+TUSG29ubdytPRHvnkcIixauEMg6dN86xop3gauRCh872vN9fJHWc
y4Azf9D02FiHmG/8z7BS9jXExHuEN2NnDVyEIVMjofbsGrDl+ph6p+trkdZPNDT3+eriVjShfum4
QhieZPvHdCHmapcXgL/9f52pI5grklex3QP4BPFhvEYH8GeM1DbDS6Rz8/3ow3+T3WV4B5DrArMl
Voq9ULIbnsO7RXciLxJE5yT2UGe1xV/a2tmwuehYAhM3/0l1vC//eSMfucXpV3gpesc16CEGbG/Y
0kLxCQDrs/qmD6zVbIazj9M4TAVGZ2HY8sakkdMAQOS9lSMBelUZ9e2SQB7orMHSkRkVcDgR1017
TG3gUoLjxtSzb8IkChzmSZGAotYSH7iT4cS2p91De1J/4FUyDZPMPl3GA69ZWBomeRVal/JfPy0d
zPpAxKH4fLP7fD8Dx99sXeAngpPbN89/Lp32tjuO9Nwd72GjE3rgtPwcYLlojydxv+CtFD6TJ5+Z
q/OJqtXHxGL6tqkEgA+OBy1rCMPYgto+f/5TWqmpe2U7mnQ2BVYUjb5sbnk7UvoWhUwruH67418t
sxI1bRjzIyD9+GwZn4vsKzSXX0xM6rlqbdRj1qEtY94ajU2J/HKhEcI+08Z/HGtcTYe/vVyRKkiz
bQ9wwzogfJBgo5+M5dYuoPP+fkM1z7M/pHb98UinoV9XZmMSTh0HkkAnphz4ogDBGh0TmLIxoSt8
0uRs6rT2np2oUevxyl2QfH1N8xfS+QhkqqwKriLocNlsBcft3XL72VnOfh/MHcKH9M99cGK5sdf5
hg+3ohmFGK4PpfhWhW+QHdPl7sKeCljvkpE1KHVVS1VukWLCizjvVNmPuGctp+0IqeN+1TfBPjWV
asJSkH3fZTvmEdL1jhSxNWcc5UefWcX79XWUBACpyikvsQu656MWUwtLAyTbKazC48GaeEZuXMV9
u3yUl/ZB6E40lZqe/NJ1atJYTpYcLEzNulFLrf4XB7rzKnOEuVd7+KBWTt0479lZyMlASEpsyAvR
4X9zxJPqOHi8N9OW201lxbYIQd6s1QuJhg+n2zBkm7VQhoF4n7Awgeg4bWGCsogQXFYa3XPnFA+4
oeKIuIXDjBl3DXJtQtiId/9WYNRJ7CKX7onBGqGkgAFdaoNysPGoM51ysjvGpPDsGAVUmynRpJda
CMPpCfzK8mQ1cWZvg8YybwrBLxPaeqIlPFEDdyI5dzz3ExfvyW3JeO6n2BS39LbZtBue7Qr2LmGB
i42xkO3OqF6XBKovIvYQgP+jh4ycYrYWMszR6NHxeYNlvTMxKtryjcymIR9SQgy6PvVqmv2Jq8Om
tagecPVbWMaNTwGVirK2JnkOUn3EPn9KIyaeiA1653a9xX9aQp+bEMo+sdeEkibAxRmj0kyub+Hu
FevTnP2+Q/pyDYb5fUDsGPwMT+DdFOtTmQUABrv1cHwCRjlvmD7bKyvy1BmQKeHgP9inO7uufVhX
9OTzpciSsilFx1Zx8sLTMq/Mf5wgeSNQ1RyVeBahIZVyExZ3ShfWjalWZG5SpdyBZcyPaAShUKsu
b+sEVZeV1C7KTJYYDAE0FaWAcXAbSy1jK03QM2/t6ylhU0TPDsBNNEZ5aBDhhtZS7RwSxpmIdb8X
d5DTqy1JQlAwRFgM63m8o2dlqXf3je90p7a50g+fOz7Djogi7wKjvh6XnDn4BHfCSfXPqAfABaYn
odXj1t8VyKZ2yH8C2UQboxJyJqpTE2E5CF8AOXbru3hnwVh/Y89ovxoy2a4elZyRkaMSpvUdyLGQ
15wlHh5JvHpVloJgKRTz7ypyoRASleTK28vAo3qDR43511zhR0OQfw4lTSBCAr7Nj5rxrJ0M4XOy
j+Tw3J2hV01h+ON9M4Bko0WrlFpGt6S1ghyss54oKji8lO4vmos0fkZlP0heZ1EuGPfRvpYcJbQo
+YRz/FFfLemqVIUzQcZvRUw1Yk0vvRXT5/DOrAFI3V36UyABLB9oqDdnP8FTykb4teXtEZa5nBmS
ruBDY64mWU3IhOGOAf4K2PQV8aziYen39Qnl6gbqeVP4Ufh2TJscRHvKj0SPimU+m516DNzPgFyH
M6Z3BE4nTA1+6bvT13YBA6Ff0AV5C/BL69gzwXjeq+azD5FmJXIj8A8lMMq98rG8XZRTcwI5yzPU
5wbByuGq7sI9latwCVo8yBz5yQYmOw/yrD5jz2kM4vnDSbWqs6XOiDsdimXeTPphZMu3jR6JzZmR
RHNcfUiOOlmRo0EYnwkFIQaiaNa452YUMBLVjtkuOQLAkgcbI2ydLxWaEQAufwmRLKeF02x4Szpi
ViWPgoZLh2ascdWl6zuzYhwHUXvPu+GdCk4Wx5MuH3nbN4YN+/fIhwj83oLDm8QrkYsdCte/+KQ7
9qLM+FrfbrekhWiOkm1Ew3HUvla/LJG5q4pgnGTweYIgQ2Qx5dCoQRGeCqIqd5G9LkYofVwk7Pyz
6pYYKNnIvYAtNcKlK4UrqfwxhYNOG0Bc6029sk91O/rkZfD5IbXFH7tEaIeOykg6KKQ1bsl4dyyr
+vfiquotNiX7aPVR3h0+lTccGCwjdtIxYFoBwslXt5Vmpiqi7CSguP6SiZcGoh+ipYlFT/dpVg/u
3jApIUvFYvlLMsR9TdxW6pFwllQB1am2I1vcQXCztMNk1hh8LtBHnV0xT7C5ftlNCwxkD+lSYAxE
1W8NIcbQyiTSpj3KoBZdiNAlE+UBxPLjy821xWpWDzvWWirUdV+UxxgoFLz2ToWM3977HifJpyGy
9EgCx7qWZC83Nx3mO7OEIVyDqzo1393ugdStntUSgRwRg6Xp/mzzusRSnQwt5KNknv2lgwWms1f8
5NOMaC4BkQWXINsZOwDvCYLYx1hMbo7NL90wLRIEVCdB6UbZdltV0VWO+UzURdqXb5YLc+DQW9+m
qzmNjiRCFBaxh4Vj12unAZrDd5p0NS/pi8Fd3tSp3i2mp2Hxh+MgkxtnLS/o4kW/Hlz9e16F+A+h
chGRAjlmlAqcfwCzIdVWuKc9ePCj1Vgc3m6BOOKdq1EgHfzhE8v8uhDuK8BhHHH1xiKEP+p/4J+i
TkbNaYqsHa80J2oVudN6ea+UjoGlj38tPZj8nLClJqO6OrOpDbW/7ZWU61k0zBn53fQtpCnjcOsp
vk+uE6sCNvFI8H5an5BYySt2vZBTYs5SKr7eGHEVGV04XxRmWgwVGSX4r9k1xIJLHyQeHtr9KiP5
pfC1VOOa+1zl5nEI3Bt1lH1tlA4ttMwM/669QY2Y2jimNoWzv6kp5zfu+Yz29jYUgVv820WkNBmf
YL5pa6Cc5X9jzmAb8Md63r6iAsNl976LJH3WoS5bVc+OjpIbYQmgvpDNcT1ClRNEimAGVYvDEkqJ
sJaOgCmI/ej00MdEED/YyJM1y3sgYM7ib4lHWwwtNrtZ/QZjxC3SVr7fQKmOKTFsZjSgCNuqSytD
JAfzmmZMVPUFQ6Wm8HaqTmyv13/TTXsgkbjk0y1uPuDm8W/doQz4+lnw1yITmKscrZ1fTCwIkhNl
yDvgcLtZncYxSP7/+57/c5Li1JzLZO236WQ8ZwxkxjJ9iiNINtwEn9il9TnxYk2TyJQFQtQ0DwQk
92by2CBnqqNp561pjJscBcXzHjsq5su/KvJtzgnQjzAiYdH/Jsis9EiEgAhOVXubW+0hGrK9vJZA
m4vDbHhb5revZPzF80qxfzKNDgu9ZvDJjVesHmPPzclsOg19f/TbGyGbILr+aMVeSLjQb0F4a7hJ
XHTqiVanGjNtI24mjcLd3MdDiDurhaqlRgdZVBzd9rEIIA+gkPiomu51jkzp3bEfviiap5SkJ/XW
P6xOWev8mUqiUGXL9WxvaBr1+UZ4x8oERtlQrguYr67fUY2ER1syEgxvs01mtZJu+Y0//twYqQr4
Otv3mFFvvgtm79PquLQt7YM6SnaJa+iGr8UCoRZCVpbbc9cAvMnPynI85vZmEJ87OGJ6zcyI2c+o
r+KNkAbq7fe/etu/eXUMKXLTxeJOut7XphuLBpJYD1jVMKDpunT5+xRos5YvxIQrtztwCdnL1Wnt
8B69ZA8i8Evyds9DAHa5CU2RepOzekch9/BbjTO4d/tbey3rZzd+j4oh/sRSEbyOSC92KiivIDQ1
TELlvhkwE1Yihfx4xIF2iOJYUAp7IU1YTYJCVyVQeEGRWrZpHyl3ejefdNGalzBxmxt1z6TeyyPv
hy2gQ3zCbmmfoscstM36umQjpYUVlmoepDYeVjIfv09lFWCiha0ID33N+lLGTE8nLNihv0j66VM4
cy64J8e7O9BnhHLIUqLCdB5uRccR7hccHKKWmotMpu34uQR6nYUhlgZM0wSbBDBZIbFCbvfdwn47
vTmVeOPymbQurpDx3WRUoi5vrCRE4WkjMkjZ+dF1455Z8dUk5fuieyaWmielVYGw2EuQDa0tmnZH
e12D2A0ogyp2/to3SSpqhKcv1IHBuYqngKEKjZzRDVSviQOS/o8R3l1shhI30nT6pUViseY2Fqck
W969ovPOYvMkCjglfPsx1NErHVt0r2dJbSv2ZNPrah63ywWAnbyCNfBHSuhe9ugp8DKu0v6UFTKF
hYje8GLAjb/t8fOPq++ynfd49AVDd3jTZmx0JWFRFznaaYO6l8/+JeK2Ybcscwmg1na2dniWcbHn
geKradE7lLDBhld5UO6uSo9NIxQ3G6hb3Vl78NZ1tb+cVruT86Ye6Wp3Q0tch0wvQqWxGHIx0IaB
fNGPaHy4b8Uqy7Lhtb2h6Gyp2og9//22XPf2buAiMpS10SQ4AHxUvcI0yqWE9CI0xb0/NlWBpm3j
FQ+2z1j99hNn5QRs2SUtimK0J0X0BCYiMJb/bhjASQDTLiyCYhmQrQ4TTbZ/NtGlDLjsaV1spgtT
e0cOdPFdExRRjOXxc72+r5cQubkSwO9zQ1cJO6T/Ofh6IUif2XsLKp8C8rtPFvwDnT3LkdCJA0uZ
BeQ4lFPDsuuYgz5vL7wvX+rlqqkZamGvrfhXe/vFJhFJA2oPMitlXNkG/H33GkJHj7IpjsNQpFW/
MkQDhYi8VYVSUiNEKPzDL/kmix5FWNEh609D5Tg38Dhf6EyM67nQfmP67ot1CakoDj+sgzjyWglA
1Bl3psFmiyWt5y1aOmSihRi2Neg7sZw3uzP5pQvoDI3zcIIbSLo7GD+Tj9+VxaZDI32icUCr+xQ5
PQZext29pNvADRwd6mwkA1L9TvuumxQdIkQBb4XGLnwL6tAtZRQ25UmGZUu8SYQSkQLsneKXEK2A
TPfdXTBLdee8xYkMzLbo5u5wWyLJWX9hqkFCvi1zFk3KJh+d8iNY7ibcJ2/T/szPRzz0ho+dI/Z5
W2dXmWsmzQG4eafwbYRIvnwvkkUBdy7WQ+Z6YnkmJhMdsdShSv1CtH+o/648+zvpLnxtJq4pcPTt
ImVYfiiFe4Z9N4mIjx5JXssznRmv57LGOjQ8FtYOg0EeNgEAWsmqSYs5Mnp2QtiK5twV4ahtQB70
kpDNyiGWKz7cuEC3HBvzfGm4vIBUQwgdFgS7/vjqp+SnDzNEu3Zvk6N0KtskehxsAWJ+71u45QRz
Etp3C6gmLsLUrnfUrPeDuv5RNlY8GLOkYkSE/E/v4o2TB1jfTnJnJ2/HuDqISq4BuWOFeQNis7ZK
NEjdG9toCDx9cFZJM2mHDY8O/yvURidGItp0Q+PblXw6YkwOA785k8wtK5ExBoEV0yQzZm3Tdzkc
yJgn2cukxz+eXSRR22gd2HWYhQBKinsXb1yuU3yvprLCVRW2kdW8E3AjEsZc/qjPJHXePMZmDMiM
xbGuTYuA0JTHqRZDcJBTvMKu0RKPuc2AHf9yGkgK+jswB3W0qNXNj4zUx0ShL5tzWjK4+Vw3PsBI
BSr8mRDgJ4oFlgEdRj2XY7LUNGMJqcxt9/3DTdXpU0ChvwCDfPwagu5uDrFcO+3XBdN8MDhKOa9l
CdncSvwU+nk+7srBlDN2ZWp6yFixEPf7Vm5JxGYcEWhN91Feof20iEGFLTl2B07EMQ2ECaiHWHKI
8Bbmxfe0qa8vkG70rOe9ipBWrYuD0glZDV9TlF4WM+mWc4n0GDeJfTi9FBss5BNMfJ9iK4Aiw7Kk
7g6uM9eoABxpAlFXEQyfBym3kVQIi1gTrf7l2xo6xydiMZAhC0rMWuobpor/VVZgwjb0QR9pfUcx
ZC/X+/OfcwqZT5S3tRksPmHfMnVYtwr6wImOFEqPRoH2Xmdr7RdZ/DDkHZAIbhQFUXeNPgmZERNp
d4g0cZQEroKL/MUDY2qtfCYx+AhNMokLLTPu54CRcRmK7AUnum8mlcDuSuYVWlLw39LqToyZOG+l
Z8n49yVh4HFtCIo03bzh9kIoDyHwpKdzpOIwHKleSah/p5U11RVUDcd91cXAXYKLlfZoEq1KKUMF
o7T5gLfGV/KqCEJZXGEaAtsBMYHMw2jtJE+/1AClcSySjCjvaMB7sNXcBIL8Bs5njLCwdSz6NBft
R5GQpPM/eNHv8XYkR7nkZ/8haXZiK0YHNMURC8TcZcYFqFYIM8iDBB9lsFKtMdKmDBKYYZf1ljec
38P3IEAUF/DJWI1JLJ9DK3zwRdTlSwfxTfXXiHuuNTPwMVswTw2JH0EMjauQivMvpD69pviT2vDZ
IHAu+M9g6Yyan9mvHL9aByrjSZEyyRpQjMufdWY/cQTaxcL/Nk7Z0FeI1vsksCUbWetGrPZgX/jw
h/fQ3t/AQPw/yQTfVLRgEJX3KB90IrlgkWLwd5AtTWCrLS0gsu49SEnlVeNIRj7cHAkGtK5NUvP0
A7QYgMjLxRUacAglhDYAx9SMlpcEzxaav+XOBCRo6wAxt+ZkRVaPt4fPRGq0qtP9F1tT9/WqXfPi
AsQ/ojDkw09FanoyhDfmER94EkCTk91xgAikTWmxT+TxQSkT9Bj7u5XU2YCsBBy5UD3YDL9hEOJ2
CkhQ+0HEuJ2YKOVM3i/uTP0t6uM3Je/9QVeL8bWiuRpBI39dl8CGXeb4zndlkTdORwQliDMCZFp6
IHns7j15Fb45/skFoT6sOlxax17XwLs0YqT9P3CaofVxWcgw9soKyszMC3YCpUC8DCXQIKuY6lrz
XYvdzCVKdnrBM6i53R928YJAILtHZHUwreAgndFEHeu4Ad3vvAAKSQwgyhEze8Mr2HVqRTzNWZFW
zIehs0RctO//achEBkVEUFv9h9csMzhEgjRoiBAmmg1GXVUMUU6BYfRIS0PmErZMyUy39MQ/jmTB
sorkgYaN6CeQ4ycX3JjifmLMr+U2xGNNZpaaUDQzxy/kkoH96LNWtEEfMnE8A+P2HwEQVZHAdDzG
f2qNC3z8RV/bI3L0TiOnaJja4v5HZUyF0Gvd4J25MU/rM84bXKMO1mGkbMchUjP1VafSnH65e62c
RfpZsNp/GAtL6CsqjL1seq93jAHFBEzWbkabsVp32T5mxU6P293VimzHSA/NllAn2gKdYxVTNGcf
FioRZqLhhaD0pdl1QLTikGsc6bWMRQhVlsNXPcZTaO5+LRyePoNla+2FZB/4AFdMnvxd3EiM6NnH
gzfsYKzIezGNM+bfiucPDOkJ/o60BprtCHtZQCWrMM8KqKG+NI9xY7gzdy38MVeEBkz7aN2Ss6Rz
TPL35HT5kkQL5E5SWxWlo8xMES6Qtih447TmGY8h7R6T0+0cn5pqSxVJUhECfCjhmDtNKJsMKbpo
lCzb9anGmZvPBHfHRaUED4A1OJT50jM+Y+AQLkrVoGZMhc91VhrVGvUNrMk/kh7gChPb34uuR/sU
FMmkvIx2K4Bo81E/mMoBB4RGTAyDRDkVz81Wb5ByPvJ5wIC1kbF2Z0IYTIRzZuOyaBGMm33KrFoO
eF6vU0mJ1R+R3ezqf0a81LpQHWYLAI4ZaBOG4K27kagEv+4SZHIaaba+TNYT9/N9yj4Rjfllq4vV
9rQCvJck5BM+pw0SrFM2X5EghR2w2dZ5Hu7VNkLtzKbeUqjh2EWDA6upLQz5UfLgLpMnmayXu4s9
SrN5xASIIkSk7Qtapd+bFjJfCUop/kpctHx5X2HwrEGPLqfon9CutYKF2d6fLlgroMHsrAiksyAS
pSo3WB47K5+enzjfflNdrBNovW1jMtmmiI1miZTVv5eGTyupvUCMjKKeDOPQ0qrsKd8rz4wO4BrY
h0BeYHd1smFNncjNDTKP6/9pCfmIKM/3DWuXQIsZuDfGBLiTC3lbhnOgjN3w6a65I5VXzP/vWtzC
qdMJ7cXsP39hlVsIALCF32yNIowfxQ9tnrkJFiYr4OM+SSUjLgwtOxrCeivgHdA2gJQpXkwt/BAP
JB/bNlGJNF7JJ3w9j3lj4D0vs1frh/wT5RyDMpdDIdzdGSGlTlkLo+xs+yoKIKiSM+3sRLOMTWxz
HV+Z0xl9d1RjKBsZ5hxQhgGS/pzqwjtRndkF+xnCxlTEqUqBY7rjM4VNErp3zs5La47u22qcso2N
Y1CjwE1JJfMqzjMkTcluihWJTW+zoDDOkkNDRESJfYsqsx+7I4/GYlSys2PErUf2oFvKzV1ZxsyC
xSQW9gFz8k0hjgyKopP7w31BpsceOuNW8Unt24CWWg9y+ffU4DEnn/Yd/AQwD+Z+TTmfvxuhzm7s
lMBpgm3c09hnoTQBKTNIbRpw3g0A66NUP3iEoj7Xj4jCUyFej8kBYqE+6p8fTYXpJu3RLib4fXak
1M84GvVjtIcIT+sX4osrvBdXFgPYmhY6VrppeuGvZrmofy60g0Pm0uTuP5eebbs/nhAYZcyUbvH7
2sqaLFuYLTOukYU92tkLRO/VudiVX8XSmvhY+RRloTjU5atRIffKmuegh9tVhzD3K7dA7faxDum/
RH5BBVp+YP9tUiQe2R9EnwT9GXSqRHG5n0BHGwKAnicBKeJY8Hwzz6pTj7UcmBq4IKTmtPvNx/r8
Wqxr15s+tqO24T7WDFg9xV8I8gU5fqMdoO0EWryxhJKUMXQa9hNPSnN2jL1qRv/4ehRlxUFz6Nru
FfV6EsHH5qNeAwJAE48EEPUizIzIXEij5rkLx1enN6j2kOsgQsxaomOKLkUoVnFzYFn7H3nOs1FK
K2WBekBTFGJVkLsJPjzb7icTosZikyDwiqlGrLdAY+9+BDB1V+FvxsMr8yoBSa4r/xJMDhANPFFo
BIEcesM3d/lLQU5HL7whwxdB00atTcHSP7CjrJgIde+oyTXQNs7OcooC4pZ9O4W1dnPkFj5EEIbR
tDJcPQ9u2keXLS1CcwjGZSLiZfTVx4aB2T1dXyszGgN8lRgqfzjbfvJHCJBTyiDLIY2V/DIFsRtK
EjKTspa8sRYjEacVjilh+eOMtkVoqVVe4oeQVP2tqRUdKh7fQTtA33mhPgz2HrovypJ7GSqxCuTn
cvrqBTlECtGVaXB3bt6BKVBv9eFzKJ8z9vwEpH+7AcaThgCmhc3dhZ3GoHdryojLxu+hCB32kLRG
NXnIMyAL4oAk9u82WgKkr7w7C4Hc0A3i6uXKjUUzGNXggkFluaqh8r4YKcdyzVA72KO+77fksv8t
zb42DEb2gzAd2o/uVClyRbyRAAiyDRGMpWURniQ7V97hnnK44rl89iN02ccykdwmppwwZkD4fxGF
sIcmhhsdx7KPIYR+GmzTr1r2n7xZQkc5GHNQsIVu/JWSxNws1jl4W5G3G29/AcHI2IfPtMT+u10V
8KR0wDnjettVPNqyYvK1vzcFnkyq+uR6XC82EHuhpxvIE97YCi2EelC03vCGxIEIHFgxf7WRy7tC
3mZC5REYIqbiwVjhgtegzIaOfNaoEfZ6FSru57Wey2xeN/qbAkP6ZfdWzfqfv8A5obbvTRypzkAP
0VOWYPGwij0m2PkLmgZdwVu4wnA4ckDmn/XLqKaFlWfW4tDqRWuN6B+1XiRmFNiiAwep9V5leB6k
U2pbM912ujfKQ5SEZ6aeUJBRUBCIPc7hZsd/Kx6+Co7eKn4Rypzo3/aCcpvLsxpTqYWqj3H89x6z
zptm9PI5qqr/HA2pei2MfZvNbrItYHuiwep7/XUB5Eqb79emwYvluUfjtfUZL1eNFQe1K2nQugk8
PsrtA+dUQCiXaem3vChigAIWY00hUHarl1s2PcnSGz3/RJy/nVc3tpH3ptdmbYnjbK3FOj8j/XsQ
0nERtczUQubt15Dg0oOkelPjGQQIVgK4ZTTIamQ4THE+f7pH0h6VBO1V5RC0bv0kbzAlOvhWX/e/
c63vBLU0d61K+26qnCSaaZeNq/TBGf5RQCPp6K+uXwE5VoU4gghsk8Q2Wl6vrKo+Akathf/GOaxU
FSRjdCyUGC78B5PtSt73QF++Dquoj/4cQw7ylYcXjaCCdlXg+Da0l6DYhnVE9T2cwZsGXEFpPLlC
zbvEgjxbp/hioTzk5JxkxyQlXPkByOywkeJo5G5qfHpGwrA+A2DLv+IqS8Uo5Wpl6iwEcfQMXFPu
7+lgVYdJbGAA6QqbSgxZVWSCYQ4uXZnzjufGOFkT38I4fxTM3U1bwkBsqYyxz8c9nnND5Umbnhne
t0d98cR2Iqd15mUzyTGtT7HWUvK9jfnO1zxpTf+s8KCnGPYpuDzwhLF8EohSuuBioQ17kwADvxob
XMDCSiXageaYW0XVbCbIrRjX8d0lAHR39SWu0gdSCQi30hnNoiTQLKWYjcoiMzCbsQar8UWdzIXl
FOygN992eFXalc9D4GY35CKuJE4rSwVpofiH5UUo8LS0KCLtfN4BSMehhf7C1lbCNFdKRVhYnUKm
YUGNCWP4+ZH5zq79weRI7YpQ7fAk8xGGcRZGOEeg1W6KPI0LBQyiYPEy+xyUXG3PdaOWAtINBXlp
WNx2uzgXT8arMRfsIwIvVfkSz/OU6tmZsYF0/u1h5XOAQohUuaCo/+DRDXN36VuJX9tZggPoePJS
ylx3QFj3S+tUegIzi2DUx93nzxT6Rn+A5kJdTzV5TCKbYAXxYfsgECaTSIyWhubWWjypIjYh8V05
xAns3LP+SBtmlkI084vor9h0WgC5lqX/cYlMAvhs38zIfoiiR5IKEtVY4/pfw7GHF2EPgldj7mjx
42/sGk4IBuZgagzn4ocrz1HpYcfnNQvqvKyZxaZZCS5mvCCvN+arPQodarE55RtiR0Yni+jppbE/
yWJmrhvdgOnJ5MmFQpjjAgizEwRkjSDUw/1k/1jX4XccnsEDhcuXdfeWbY72spoy+cXU9UHPIekt
Gt2ejYVuufKENhcS9fYc4FsRAFahe1g6vVvPBU571LdUgCjyObb6tktyARXD4d5aQ300yaGVzHxW
QTWqcslYp7EywyGjVZJ3cIXLehtEuMEs/jpCP0DcGAoAKIjujh3KNJNu+p74/yNWf5i9ylvJ/K6T
71enCTx/l+HZdI/nKR7tHu6QKYloMtDvX35/Q7RT/X9r08NssSo+weDC8+bZoRqnqmcwctsrcG8Z
uaedkKc5IfHaOno2fwud6aJQIdUo/cTRmxYC6NBkfvbEZn0tf5/em2FYdcZepetNHn7pjoZdNQ6N
wfE5XD6+OKrMte7Os3/IX7WyRG2fIsAOL0ENcZUBtiKGNelKdjPMZbWVYd3xW2Rai9EtQlja4W/K
Xm1ghdzk/Uz1mjzrC6a1cyfutdDXZtZ3hFWthZCkri44x+U7S5e6tQXsRRHeNNErOIviL+8Akqs8
OiALX8x6eil6arKhu3RnqX0wHZRVObxAPFPTG2iTKluuDHcmfwLlrIKOD9EUE9gyVNc5YOndG1iT
9+C86Fltxw1D+IxAzNlbUe9JApgvmXZJu95OIzouO5i49wan6RRIvFWG0+BmcTC1CtA2UlTScQPY
wSzEttwA1o0dcC7A6Lw6MulDHKed9NV+c6T99PENHb/uaU8eJRztldLFBVsHAq0NrqYKzoBRGDBE
47libT8TDTCsCzv9MYJl//XV0gvvRCrKjKcs08CLTpYQN4BOZG84C49/RVMOo1IVoTc3cin9us1s
uMpi+tXfKv4DgOpfCrXuDuXVyISk/cFfizY/JDv9NpQmr1cVPz7dnROC/YJe2LaJR5R8KS9ej16T
kO65ynV7byvQCG9zBHCWz/HMozclCX1e6IzoSZxoXXL+ZxJCJUwJ5J/O9Xd+DO/gFUUo3n3gzwLi
K4G8hrsrBfVzLheA/Vhx0D4XEgvh/ex+RTcfBxDMtwv+40lBdEIsjPMtk47cZ+PSRA0z07kJXWCU
EAkbPg/LPfsaovDr6HJfGYYAZOvTtVOP/3PGPgbuu6lIRZIwG+UrJw/dWsbn+Hpf8s4+5A2NsOet
TI9PWhA0PXZ+ObaIzbZN0yBuzoAV9MT4zSskHmQ0sgX4LyiHWeVU3mx4ZnUYWJJdCkmCdJFqo5P6
9+FMG7WwDWOYaAoDNClXNtLaEAopsng8Pf88dI9QcX9YVwrJuQRzqwJNb9I8EE5fqULCM1BkwjRb
6zIF9C3p4Jl8NiKDiKyCI1cy5o2BFTjrMeQO+b8/eTF9ZugnGAt3G3lYwg6oMiyjTTDdw0d+XUtK
YtPlWn0/d19Zy81eFDWm8y6+QpVE5I5ncrUpns4oa/+I6lOwXJxgKhAQ5fkFCOug+/2p2k1/WAzg
XMCyciAm+fbW4OAw3ruXn3W3PZPifmHlJq8eFqzP/QUOXKo41FdcMg05cOQaDzvOPzpcSioXgAcs
N3avBGtOGtR3y/yzsc7PFCGTkcdWT+2M3qROAA0N1IRdqdLtKNalbnrPOI6OLYm7pp6uZuXc805U
r81i0pez92FH5fT2+Q8W4NTDg6LrhMselgP4Z1LNeIFgTnNtSp5Tw2AAxi1/Q0o24RJqK7dZ7SVL
yTkZVAxhIPfofxWZRuDkeNJXpPwVwGB1xAqU47k3mM4sZDEVZcU7Uk9C6Q+GuOiGfdVsSxIq3dd7
OdfNWjdTgq9oQJ6AYmJl7nNrdCtZ6eAYlRLSmxTDaHz9/VgbONdEI8TVKKNDNMiVD+jTvLbkpNRw
uKrd7c2Nlt1Kk1avm7MdXMcPpdBCteIyUgtkzpyMSz5l854vO6k7sLsEP+Lz1uZLrnirgEXaybJJ
icoc+FUqcwOmxcCIsXJROp3VSD30D8IrDOo0daQ4FGQEv5ARU52Yo2Fn00Sd1PpLkLFBfH+26zxE
bpr+mnsgp6mEsA61kXJPVEPWQogJFbqk8/r53AY10AziqVKH2J1Tbj6518B4srF6ah0DQzNONnLg
G6q9UfECoO9t30M0NgkDqGuSqJ6LE5G4kgLlHCD5V5cH/zmkoW5b1v6TsSloo24SdmrssPLAwysJ
DeTFGMrw6kQQ9q5PP2ym35s/1OnlmLgvQV5s0KV63/XQNz1zrxhoOFB5eNYVBbMkEDfVRbPrj32E
0DZY/BOu/2tR6ACZfott5svzasVk94eXd87U2jKzKuKrqtnpcCoLsqu+lKrl9sAKm1xcbaabFKLd
65lcQCUyJ3Fm8ulNGuUPUaL5XrlmixqDNGJ++2w4tMrWka23E5wERDVQ1eFHrX4U8Rs3MYDGlzHr
I3/3LeGSR47XnOqV/ejAaV/SJfGFofwiRiaHUKjbGXTHtL6QHhFix1vOdOvHaMbU0eoX8td9Q8YA
U8fZbeoLnA24eaPzAm/hScht6g/Uc6iG1JZkg4eOoSluD5vSvGdxRjWEDvO8pGX3RwdQ6LPW+5Bl
dJhd6u9uDy0qIHkHG0O+IE5vrvwAsn2dz3k8T3JKAmWM0AX/4+Fib4Fjl5QdAON/fBc3BuQ5oJAu
raHfrXcqQuQI39XzEn4P51Cm7beH22pws0bFnVlDTcy0XCKDHZyVYu1h2J16PKL2ZpTU6tXtJNxR
hHVFdtC3+IUpQB87puRaiDAUI5m2Jcy5Quy1E7FhasJDk8qQclGxOy5NsZXVCOH14ZJpd+sZF9Zl
mRlRSwfCIl/A574MzEh+I8ef+WCvjSWMXDfGxM9h1H5aFp1a7QW8iGLIv7yPVHWST0il0pgjM/2q
1iYgXaBNlxyasjqNnnG2195GUDpRBq8nYHapK9OUDRQZasIAJeb0As0c3n2Lc1tdnyPaQQsda1QI
W0CR4u3F4UR1xNQ5UPN4yk23v8gnHb5Cz/7fDL9KOzlvuEZ+z7lVNs2I7kXuvTWPKTg+wnT+PETL
z4QSlq6npFtra9M1IrDavCnXFI6yyq4Lv/KX0BF+rfiEmqnrMwyFiEW7ENfCbifHagIURNR8Ls/r
vak67yJGIgF3XB7ywTEeQMh8vQB67cg7avTedCH9a7Up1BfwCTYFLmRuIulWajlcxt5EKadWS9es
zBHBevQntwtzj1dKyXwNaNZlcJds4pBMsFB0WVpylbQ9jZ3lYImWKMfNvRiNm7/MDthXYHVvTfqq
m2noKnheRYh95TJ50VeNUWlIxvCknf88M9smu2baH5dMJDu4rZZxUuMh6v/QDE0K3+nZaYLSBzZx
OZmBbT/zoxFAo/IPY2oxBn9aXaH84pu9aq5c97tFxd93uxSWfk2euoI/Bq1v3+kWM/MzP/vL6AeQ
AIWQsxUzHOrHhHIxvuCit+Hh2GjdRt+u7x0OFlyb7H7UOON5nXLm2yqoGIyUD3byJsLrvwqVz9/k
7BAOmPjNw5qzbhMO7vR5XEIjMUBeoDIi5kyH4TjPndzo0nhJFgxWTYGES0b9biNB7jIOTPHuKQtf
bQXgUSKfqIe74mFvznRU06yBABZFYc0lOdiOhsBy4Gft+TVrRVQ5gF/NGjqIUTLN2/Om3NYpTGT1
Dh1fcjX9HRD22mHSkdMMVuZmC/3NJ3wx+29wDFu1H1BtOndiP0M0Wn6b0cnyz3rR245Mw8mwyytN
c7yXibSBh2K1Uvb8ncD5jJnbWHo1zLqKTbnDxOfr4FDIo7KcFrpYr05Xrpc2IXi9twBf5wt+Yl10
PaGQd1dj7ZvDAUPX6lOZDWq/COZaRfmTIOzYMAzr0fi/a+lruDgm1THjJyMxPAxKICZ2Mpt0Xjfv
Q28EBn+Bia3pGFT2I9FzGQ6nFqUzFMLopmd5LvsSemdP1PPeszJpJKPMq6PdnlBtWolqtmMHPGXf
hDxTto5AiMZgkwR4xj25+g4nFIlrp3tCAJnapkpQr3ZjMJEpCeQP8WaB6XkeAGfbVzVQ/hK6Qtb9
fyegULjRBjhM4hHGsfi2WTkPqP+kspdACc2Wk5MFzktOhES7pJSe2MMwGmarVMaF41QAV7H/gyOK
UjJy2qGywjhCL9nB1Eeii++k0qaXUwFR6A3iEQumu3l6k1KlgJYBRON1IulHVWmhmFoSeo2H+FFS
Hki2Hvopap6YEDb1B12ElvqQtCWoZJKg7yE5SJAvqgVIpgkbQyQtYxXifxA/5dUWWMK4OI08sDtF
p0I89Az6VExqEngtO8Aa6xOTbRzhYswua1ltbu2Ze0EKEpAhKC54MdfeaIvNSM2B4z2OYqck1Zy/
eQIgiLo9FhLyzlSQYK6SSS3zmN4QjaS8Qa+z+YuI4K4Gd3C3F53RgBATPxGy/h+ftv8GwdCWpyJl
7UFUhRJ47z7a0J3DJd8RUhle6tfMmtVDuPOGJii7P7RcDj3NTU1eqtSFmRDu01rP5nhwBV4AwT5T
Ejzt1h2QCGJ05L2jz9e2py813TT0KQJ6lSiIAdxkI79rxmAIElMF7AmwdPg01p2uG5PU3fRU8442
DoBmyyGHw4CqoTHv6W8O/tEbcwF0t4Luu1k+nPhoIGt2Gy0T8E85c1xdoS946tNoi6d1nwIDWjI8
p9ImBRoiKaOBASrMvqLFAifvAq4vHl5Crfd8V1HNEhR5vEkwxglyTaRaId7LDblvY2ouyyQV3O4X
HhF1nFpV3fNdb6hksBbj/d8e6Fm/pedYT+st69GpHykbtaaO/6d8aTWd6kLy4l3CJ4hGB/KARiFq
FjfVcS6R101WtXRl+uOSs3Y4u8yUb/lxRplVfkAE75/DBXEJZDEydygU4U13JufWO1QQR6RKf9gf
81qjKOSbVZSc5x33DKPhIM/YB+/AlnHD085XrMpUv6UVzgyte9ocGREj8RpO0vyOROkPfHUYknG9
4dqjqsLxE/ZkKNcB2HbpmWPcmoeB45fr4NmvxRVEAjPE3JrM5+PNrjIcRsHEEBJ9ZqwSwfU5urG2
ruuzTR/iL50HG7rSxRbG2X5FfZ2J2XuHOPknvI5Gyx4xbVvy01APPgFQBwGj1Vhb1NBD7/x/dBM8
1WrXCvKC0hd8MTRirFjyXMaHh8HAn3cDa/bOf09mU+4U3O3qKLjYT0jzy1K8cvxJolLQ6M0CUs8h
sgh86IRXnNonIhHhtyCnvcoCfMVQWY6MchBgUIZr+izEFJ3MJmL3K7TgJpkTfOhfCLybaPGH8Jsh
G6tg6HvgZJiwAHyVqfF6CX5RycDGijry8tKJy20RtBZCzkf2YV8sCdzcMzdBz5UWIlvBLxyBfZa4
T121S8KDgdxsqPHzPF+dRJHwYHwxcaDHtX0qGDyqlwi1WVBIK1nCGEKUUQU/iZVYpNqgmOgZ3qq+
JS3TFLMg459l9WCTIny28/pOYm5MBC4o5plZK0aKQvIchCeawH5kLN1GU2UJ+RW0YvN0USRD/jQ6
O+esELxo35vqhcET/C4sJvNwWzcvtgpyAHZflt1H1ARgTu4gDI3i85Ukt1IHWI09Vf16g/HuWrwb
k61JYaRV8r/9wD03LLJFLzLGWau7RAEmIHBGm71YNDWaBn3YiPNv1LcvC/66YsvGpn1rXVkdDk8C
omWVZhvM1y3dM+UHABYJKgj1T39+Y9aN8U3LLFtoqv1J7V1ENisnJ3gnVYlQ6rf2gdl68jaZrdiP
AdyudxJXDofbTBqqn29aSuPMhX/nw7HqkXtn3v6by7tzswN0hMgEWulKGsuZS9UkfAW08XLaFGq3
ZVwd+T83EbghnaNVZRr41wSWUrUY+lHK+vpM3H25yy/ljt6se7VaULSLaCVoRq0V8o/1uBWxfYLI
PTH5j19NJvb3xxKRCHmcC6VyK5jDUNskO9VCuJsj1hqbQEu2/wkIwf5875iZ9cb3WZeHZTk7XkDQ
wk34lVVWTLoTUAV+MMBDVgsB11t3fFInsDnLmvxN8l7IlITOI0UQbfPpkTcGE8UqttxS6/u7FyQR
HORdmL7U6UQXjaUp22jDjBh9N7kPRVRtiwnXDt/wpVQ38gW7mZ8oAkp3ANZ8h9q1Z88J5XfuU7sD
oPhW/37Qb1AxChNbgAAbgj6tmkydumlafJybzMdIUqP0xTrZ9qYuibN4k1vO68d4NjOG80PXtWUE
GOnBr6brldw7I8Q0yKA+ExZjif8Xf6P5cvDxurEtKc+545cPmY+lccjIE8dqkxKo2lTOS6TGgJ2n
87x/jsJSKesofb8be5/60jtUh3tWT/uKAbOcilTxXyC70QmUZtXRujC9JfQZDClRV1CYiQtlkfAu
WP7ufyLn+Cx+UAsCGpKhzbVz1XHar5JzN0K2eBG5zE3j15QOhjMRr4bOJ2WNVZ2nNvZqd+xyxKkb
PEJ9ZempUqgJydhfOKVNKKq5MkBs5fLeSH0L3xnnkc+WI6is654RE7Hl+f8yPsxr37BQJOiSmG8/
RgMkZBu8pr/HuuudePlfhhHSmTQvqJliOhxDUC5nBN42FLzfhm8P80dK7BXlm6hPvnVQ9SUKIE0z
K6/Ee8VesWF1tFeZt6kTvopPqAZTMR7RC6YhC7cs29xp2U6xm/yzWZMFFSHQaC8Xnjgxiwf/Ws7G
dbrgYQ54LDVm7cvciLAyWqJSqLUQwJlK9ev8ZkWtZz1Ej41hJC5IFemeo33I+j+5f2I+kN/491Na
zXtv4e9E5N00PcGVeAZzgxyKGM6R3Vb+JBqrAJIWr/7oPjCkzhxUsRUjGmb9PhyJKCdIUOS9bBDe
+k1PvYYDT6yP6i/a4zMhTK2ImhzOoiKB21BcMlV4GmoIMj/7L7HdWi/nAJfwEaRLp1eHib3Y4/D0
iCEHn28ZNtWHXQ7p5zu/JxoBjqO9YTSQZHwNGAxuwpsqR++/jZl+4xssRzxdzdE2EZBDdmoNXUtR
NoO8ScttYYbJyX3oVjroUR8g51+KOkMwYIGdTaMrGVkL4ZyHOeUpalg3rK3r+RDNpeWGqX6G22zS
gzr51qlRN9T6tFr81qXFKsDuBloDJROwrGPDS+YCWJ8UVeiegyjsm7ncJp+2Y/8NesnCwXJXfZjH
W6ezDIchqtDsI6wRuc8Y/lIbP6+VSdhlP2mIXg+G/lcqOGuhGM2Fp7HtBuhpdLRgrkZDh8dbTh3d
2EhMdN5xQXxO00eCZ+8gIfbTAKAFlSmIEwX4s602VkZODq+Wfvl85oTsS0wSMgxHqWiOsj6qHray
ekn6nnd7wc5I1phx4AFBqzEiyrf78ok8QP8LfIT1padJmDWVnIQ7AVdzL2yvmlWrfIjP6YFqLKCq
4WYIrgTTjUFwMFC7WG4rJJ4rokhb6IZA5y4OSBLJKMg/qJpPJpGBY0o+9YvvXEVZzgD8TK3BO3wl
KpHqu/OOjkeOXlUUI5rV7ZL9hVMkJegDoDPEVcCYFdPYWb16sk7B9a1Ox0oKCIuSIt6cXazfwFkn
mSHqN8qO7x3UDXd8oae36U7ebYu3p4T6lGbkmu1z6k77NgMi2Z6liHfOajoTYRLu+Iwu9ta6CRYn
xF+4+K++Cp5KPoLlbwSV2VjuWWoQYw1KmhPreMynAAmQYNgjTNDoW9oc9NxAAEa+58+G2VU+1iXq
4gP0+l7LOlgj1L7GMBCXi1EuFlfNyTUDCNbnJmQun5L2o3BpYwxpAVQxDOLvChkIK/UCGo/rQMPo
TPz+GSUoX2vMaxF/gVYMQnsbT/qbU2I4HnNqQ+PQVyDs+STuwrgyVR5C8aS7w7SPx7wX2JwgwLRw
v1ouVeLKGhH3/sVo+6kbbKL4p3kqYyAE7Xsz9UVxRTEc3SB6EMuTRsGSQsQXqgq9cktnw49svjIQ
s1SuvlQ1Ex+PaIaBcC6Ksbx2PjoZ0XoPZGR4MskPQXrUYYnVCjBUisFMGDlMeXbXDo8FAhfU6Kej
KDl1eNt0XIiJpvCs5mtVPJ4oQABJOhWBQpRiZl0XhmykUB8F9q8tBYlcbsSrR6HWChIiiEekJFWn
jnDjD7q1tLs3ix1Vy1ZYyT/8UTqoxr5wPINDQgvXh/cL+eOSEk3uQ1Gi590mR1U2A539ezHEqN8/
aaUY369zBv/coCMf0Nk6oaXOaNi2lgEWkjlbbADdZme7w7djJl6HkTNY9+riCJeCWKGzqPzDlWQo
Xz4/p/OK7UbKAiE4EpjwunLjnzQur/XVHm27F6olmgz5FeadUYmn9WT+Yp6OKhCreaBp/ZJt6FMf
LaXN7E4ajPspwNQ8Pmlh9TNXfkq36db1WBoZgvqgq5Ga/2AJfvg3Rux66GDAyLBafSN9vPh+dg3J
FMYerlYqvAX2UrWnNmO0oR3gtMA0ZjivYXAb7djfYtc0cUmQGx4cydQ4NBUFF/SKX+uWbo+W+sQ9
sSq3OWO1kSe3A8/Fs6UcK80NLh/iZU2U0VmlqlzLA+dDOBp5d1sope1FO7SLyVnSPOuS4u+vttWe
2/2oQ/MdYT+srRrZtS/AZN8M52sdOkwY2FmH1H7v2QCsKLZcH6eZCwa6F1YsS4VV6I8WNgGNEx+f
poQht0l1z2HYl3JaPtzOMvlG2axpY21Wt/LQqGNW4jOcrat06PynF0j+kSPqyLTuK3iWXZyOs4WU
27xgtV5085dvzUp+yajOM1+9DOUtg6Xqwo1D4g5yVO2xQLftOQjNBJUUq/e3qxbwEM7TrQUI2f5a
oAa3x6xWMRqgNqQId4uIcVhVhzqH8w/GlNAKmzjDGJIJVAK9a53YDr0ubSH3ALmXiQApJICR5WHH
Q9fIKfv2SdJsUgg2YQRI5OmCbh9csmA47YM6F1CYfbRO1oxuZqmtc5qU50xmZQyRMLUeVzKYnQ9u
j9ZHX94hmz4ygfwYzzKXik/jDmO5PBwBHyrxMVCivonE8krz5JTyBpQkQAdJyyM7UYRD/KK2dkVH
t0mYzlkIfIEhcBNzZTvCWSAl2Rh4yj6txuI45GYCOHCqGGL0UzHDC/gFlNRnTIzq6eaMZ+ZcNdlM
OMyhGTwptcAcyDStOb+F17v+u2l02ZNhFP12OrvE4wBLzYk440qoG23SxwBRFZ4pK8KuanbIOCNf
HDpw8Zrd7gYAMMQsfqRtgW2Y6rrlthgxWoo3FVrQ1LLYDJw6YN/TIlS+V1XrW4NMyEDxCAbllO7L
TYZ86ySK1M4kAR6Ft4nh6ZUJlbT3aFDTUWBF9EA/XVAVJrf9dDtAtdQ9axJMBRnskVjD60Kauled
CRB5l2BWnlKh5B+NTk9aVzgARjAIWr3nZ9Z/cw+v+7mbOIbt0UOkQ9wjO2EZe5eETGSMhFT0B8It
KcP8IJ74/DGEOYLbDZHYsqZSe1NnccPcB6bHjvnRw8hOoeRXPzSupjunMJpV6acwj/CWOy3pgsS2
d5yb2LmRt7H2u7u2mYdQDPy6Y7IkNq7kJHTGN93maq7dzS8VEehNQwt8IDMtQdTBh56NS/R5r0/I
BJaxco+Eaq1oDqRGV8tTS848le9KEBCS/tRYFZlvnMpn2YxJw2VcaSbB9qj8nsofZIkP19dEB9iQ
hKlo5i8jMLmxqv/3zs4c7qenATVAGYL5+xHkpoFbn5OygPOQ78RoOOA2oKwWkiOx7YjlE0EgXAlg
qO70+wZzjPzORh4UN1YdPyGHm4e2XTt7vHsq0DBvIuTKYdSYrr2kn86YhF2W8AbpRZ34klrQA/Fo
JM1/btQcwjiX3lWXSsReBRlJJexq3QW2vICtSLF9/8hR1NIbqSwQlbrHbKO/btM7Ki19VO38jDtV
msxruk8pbnIH3Goq15wc95Qy7Lz8HaAFhxMQCzLzmAR1srQPlYupZf5aaPMXwmKastZ5k3jrLD2H
vtE0j4kaz7Ip7OnujaYLOwrSEBk2dBIzqqPoLD7TV/YWMxLl3P7uZLyUGcmX4bT9yuoPW6ZhqbKh
43lYDULB4cXID2yXKelJyYF9uYGVNVRO/014WnSq72EpYV3tnCx9CFY8pL0sw2cSMkUGPQmhu07q
/tUbhHHw95B75xuqlc26EKIjNpITlzf3eIaN9Q4ubYTJlN1sLSuBUWD6eTvOY3qdWw3PKPuzxiMm
3sTDz9zo1UA8qrflFXNYfr4XzafVtK+l6B5ygB67c6Pqy0MBQauMZBdX2V+4h6966VGRjtJTX6JV
Yj3rCl9Qa6qNVwEaWMiapIrZK3WpylwxS9yVRQsLvUfFjVVx8+NMOHu3j0rbJ9CQdEqvoxbh97Q1
W1RuC9OXVKdrv/D1t111zSQ8ia0XAPtOpAwbw+wXdq/Qgu7XJzbzvPFrLCUaJiWsj4iGitVtz6D1
gNUJbK6akWyM6J/zmp8CXoqF79eDlDEMQQqXluEQF0r1Ho4Ua/LMzeFYIhpRcXXETNcAfBlDAMq4
xC4Pzb+me3B0dVuZmdj4qmTecfOv2aS8LYQeSa/kAQ3VqY18JcMc4kup9lJyhLiMNnZd9bJMk9KY
fXmjnRc+aQ01XIqxbsgNaoerBUsV8Bi1xw+GFUJ4irVQPk6wOhLYzgkZHz4jKLYima3IdxzwnDoj
pZcoPOWRl2Yy9YaiB4E3nQDLinFS13csoHld7LOQjG/a3pL7mDIo7WnN65YBEmXDMVXzrz5ZxCwh
0Rcaez8BxVxemuCe9X37aXHIN4qdf4A3V/d6gxV99l15JwTPIswzaXdKte9109TZUVzEwlgJwH2J
fiO4rhGAp+OBws9JASsZT7k9GT1MELX6cB3DJS+0iyyreuyjlYezlYJvTmSChXGTsntShei+WE/R
QDcWurQFZc30TQlLrOEaZlcWuP6RZ42CbETLm5j/wGIH8XfUnd6KmBjPeJvzyAKQi5K1wOj/PHiE
+spCoEfMfhd5Bn5RZ75XgMsS9sWvNcEP3GKFKlCzbmeCy6Vs0pRjcy2zpE5/zHkzmMbI2Ofog5g5
XqPoS7OfZxjlVBk5IpuSRuLUD+YmaKDvKG2XG0nT/iBmY0Loyek21X3WwfPkH+rI/S4/UKY47DY1
X11wQuI8fLi8kOdCHJljOSatDdzDQfZvku5iruauM7XRFcgw5otDIQ5qN2E2SevGk5tXaOg3Dmo/
peNuDxCnP0FGHhI3mDyP0urIbeY7uWImY3q2V5QhoDfdEbSmFZ9ZJQsDd8NNjR5Oy5m+bYh+d6kL
8ugmFgpmqtvpUtKLVha5BQkUsqtTfGmh0TDHkKKAvoxk8etjVJvmbKAAS6GKW/RjY4fnwt2P+Gna
2HIfG/dMQsELheyDEUgYBEL18nrlRx2J3nE9VaLfgqiJ8KHdsyHy4TL8zLGdDcbNcPq0/JPQ2zZD
7+sjlRuEBTuwYuf9Pxu+AlibNNzQ9zEqp5IFdSX2KDOjqb91dXdrK+Tugfe+qdANxlAleaqNpBdn
mADtnw6M2BpRoMZIfCKk68NNhqZvnHv4VxyMlvYDeru2lvaR43+mqPBIo4GqQfBucKX4ebqigvEr
GdaT3WK9HRGRu6+J2S7/tUU+YtoNidiNIloAHpva3Q1vYy/Z33UR4kYyc/UgWhSkAq1UwEZmHWg1
G2QnzQKNlKASR9vWNWWQoCwrZEFVPPfTqVz+uSELB/me0icOHJY16OUXMdO8o0wmlUNyFY5GpU3/
ywOD4Y1Zu7pa4ddttQhMUBQEDLBHuQqUHgfLf65VLiDmImdxfHmtZBjACZWTEr6UuOfujfOv/nEj
+W9fU9nvS3c2b7XhB+Xq7NilbMfxzO4GHoDQAlOHkSEahrgGadgdW1ogJUrE4FrXtcSIHmXMO8OF
VJNGAs29XesTQAxa/ZvybWQaJGndvrAmE1kN9EauuUq1dCFP/3OVskJbBFobttHha79aau0fXo09
goSGb2TjUocE5S/sKsXIxqrujE9vzbP3WEApzxqKgFJ/AGIdWefZOMebvh9JpVWw2ayI/XAM/EC8
0RiT0aSZEnBfTNTy0pMur2LYxRDFK5CUKtfPDIad5e3LCtDkytESbMkLbw7wlbolK+ho1q7au802
V7wKL3kFbNW1sLyiFLPw93zU/M6F9vs4u85R6DhYacv/MJNL1Vsc1yIW8Ugfm5BhTYm5CgkDO28x
jbmC8OOETO+k13ZWcp2dy/UDijTshowHSpaHzgKOLYXZTrkKpZv5YptFdSFqSf4mqFZ6UeLJRc04
fVTqw9MaxzGS+mj2CtP/6ywnqv7Qb6Uyk9tTZf9j8bBBw6vJocAfn+enD8YOgvm2ozX8BryVtGDP
iS4/aT7ZFvN+WdDEb25QjCFZ4hOWjVBRb5VNaSpKd1uFUu05nrDf6YxQVZyQluydvpEtWi/iuiFp
eiQ19qzFBpELY6Rr61lN2HIIlmO1KUPZLagf4zSceCtzCP09D6p8eef6OsjQOQtyC88wTbW6sQQM
l2Do699t5w9K6eahL2isjzi2xCpS6K0ugmKO7t+a77aM8Kgdi3V6lZhs8CfxNPkpEnuyxipirZ1n
7ul4hln/5nQgg/sdjh2tukZh8HE6HOe+zLi3zaMdTsjHrUX8pBUNS4QflGt1ZHHbDktWC5uGSmNz
beNO+HeFO0zJ40SpF108aGtlwXU7gY1L1spmaZfuDK5mRwcEPOu2LWoL8ciDxF8G3dBpeToj6+uy
xvGx2blGji1h1ZSeJJ783RP8/l9hdQaZKmiHwzaiCii+krv0d4pUPLM1h2Ev7MklM82lV+oR963c
p/IpHH7EVl4R8n1mfRexi924/BRbB+/mH9+4gXxmvB0LKjedOdqYe6xSerB2nsnrsXSmvQEEOpoJ
deUT6SzRzFV1pw2EpkOcflAQDyE2YyegGM5Y+CTcz6AYjjWxIXYixPK9quxYUAglWXZYEwtmX2M8
BiGQrZ0PxnPWj7g3csIqqrtBHPnIfJQsqLAq4E3MYr4VBByHfMsiGDDDvM++nq/vZEambwxKKrej
NxQCwXeCkLVhE0Hl3bU0xvtSvroGaw++VJBuazcbz0+u5y5LBFz8bq5Ecn6DfbgtH8pV8fEXiWdC
hUOFuHzei6gHd2cTQ8+EW4RFr0d4J3ghbweE7/xDiqt1gKASBVbawxCy7dSUjo98myf2F8dZvjn6
0wdUrUqq+irFCe4b420v8vqikTRsqdj2/SJp3QQKQgYL4YYaOD/KPsY3cUj4qBuqMenCQGlm1uw5
pR6S1TPMeBCTHWRDXWze4BY2N56l/Hi0/tGY/P4D8C7Qk98GZUBQ6Vysry7+F7U4XI1GKv0g1f5e
tGEYqthmDu7I7aaC3PhWeQGzfxP+AJwdzpO3cXoH7JwhXCgvEwEO9QsBaKULDqrA177YQQ/uIqrS
/8DQpXwCWdAqjdRI6CDgeHT8CdCUA29AD76PvHFyHE9fmmv8b1ZK4BpplQ0ke5GOZ8OpWGptvmQv
BCmlwquUcYvU1zFkC5p9VI1fw17vB0fMGT/nsNda/Kb25EUleY7THnpAwuPutGuHVW/wR4Ckzt/n
IHUbKkGN9829y+GWfoE+sXcUtjmzHdNx0rTZQoLRgi/WzzGI0diGZBFyBopKcQBj7M5AXCO0QRmu
w0fOmjnv1NHKJQQtHR2unvkbsrmkAA4VcplFtCr464jdK6UDJQ448SqeAsfq91vNn8YQ8atOcRb8
vWKIHkB2r4vAmb8OrHlchqFjj8+ttR/pSYM3lLf6V/J0UnTLyoXDqBwz3dydFYWQBb+rDnJgIyHt
xE4Xs5EdHTnskPwprhoXEq+V0wQKdMXN8iMmKXhOm2n0s+e670xXqmU+ej99LNmh5LXIUVmQD0V1
QnKdjyS7IEKxISdQtnTMyDt4aziopbpQIGeD0P8SYF4qYY4NTEp4ceOuKByR+xokNucDXIOYUF55
Fh2ztjAiU++MIvZxKdeqiSZUjNZxeX/wtmdZwY6ntc0CKQfsW6ZbTsqMYmOdMr/lL4Nl6d4deJ6b
k9TVOC5sgXzrsCfv1nWg/j3O7SdPvxoSjV1u/gBQnwp8VR8wyVwYMkSUPiH/k2qzjJHid8AHdwR5
aZfpmS9osihBwIeUH8dDKL1MnBPuhHhy+l2L22qQvCBabLSogMp72TB0QSPC4QYb3dSwQToy/LJi
WZ9hX/UB0Xy3OJeieNg3YFmxUi9EaAyEpZxz3RmGnNOnX54IPXngr1zV2q9LdYSl6Wd8SyDue7xN
w9wJu0YS0eLzz4hoDI4YXe6kalyPfek+PxZ66momYKA7BaJsefPf+eXmgFW0XB7sB0vc0fW2E13q
4lUG9/vZWNqYnjSDHLdkI9f0z4uRvPKfvx1KPYuL9XzeBc2eTFcbPZDgjmZ8c6HrsMULNVhezt16
7eb7bXNS08B/0z/7RozG5F3v5NCZKQTNldqVTAPf21IE7RRZsuIwt7jAT9GbrmK/2AgJz/8kqNZX
dwol3xtoMQZ/AIyfMf6ITSSyH5oKqC2NZlUItqVW0sR2APvUGQGIeJmH7V3efsfoK5HmW+x6dHWE
wtkAZlssq8fEEg8nZT81umZng4yJaoO7tPyBxS2T8xjoXRsPLklNrFsS+u1wKP53ESb+iedMuH4M
bxNMmulrwFPAEoKSl4Y4amKA0C4tJHKBPrwFvHaCChhpH0Ay5akMd4ZnU5V0pPt7TK3HN25vzABK
Uyz85gB5SKcTdE2+PovAtvAU1K41RVAjCw713J1G0/akKpSJV3yCPOxBwshRlZwbPtipUHAJ5TQf
/cXc78dVVXeE91EtC03JPS0DRpUW0YM1LRWn8toYpnwg1gsv8FwS08a9bgH0m2hhHGaxKLww+KFc
w9UpOdd4DhjJdB/NAFdegpkmTSY6Kboq8fvpUYv0XybFaAYWERm7QgRQOae7NDt+lSroLrazh3RA
W3aL5CgKQCbb3IZwSw4NCU2ATnngh///GXh80dh+GyKBi88rBh5K0Gm5K2gm4ZkIQ+9WCusIcBwX
DRuX/tPbU2ByN7uZcWyBD0fNhObki6Aqmr5eGWIRKo158i6twNu12L9HGMsYRIhgSNxQrt2bOySP
6XIsH7WzvIADSJfdLec1Ze/S7GTJh6s0G47NmXoRRbOY19tzpeSiVs42DwaASLXZGNEb/sUZGAgD
TKPRUcEgcf7voJVWfIRp8h6ySOiQIHL8s3hoslKb6d1inUmMRv0ouWFPH8avN5x7hnPa0sQIlsqO
r3xcOvxehDDn4T3Acx3rotXcpOyjEJvIPiD67Mfam0cX1PZjprEkiVRddAudM05ToHDXpbyL1gAM
LIynxIErI5vKsielgmSGDW08NR4m5a/5+hFejmsLXxDjeLdUoMHootO0jkZZXsm9DUEMigfja/b0
h7+QspfJcdF36uQCselST9IVJ+lX7xD6KPx3kZMJERhO/htDCtgcErdWg+3cDkIdtYt9YcjL7xPg
vk1CEsz4+/zNfGq9R6DlECMOGwi2AATBMUXRlhqCa1hysVZzrM6SyUsdJjltmpXaKfyS6tacXojz
P1C41vAJTVDI46LjA1XzSsjQDPWT+r2N5+4h2IIu5ezcYVWBXG1DXF4VuZoc8eCSG7aBPuFX4/IP
hOYjGTR4RJfTrJBbYNiZMOSz7VIL4rulD2V664UjTWIpaX/OgeaYxo/gtphcnAIR5Jzr1S1RkuI2
TCd4BsPGjSdTe4vtMpjozbUpQklYpiY2Vn9CO9q+r5NxwxrEqxZQcHgU2nSCSMsjvBR9+zkWBbjq
+o5S+eRb7u8DN6M7fz68d4Np0MwuHl08LTYx/asF3WdoTtb7Mr+ygqUV6Pts/toVtFJkwmUyX+H8
tpxzNLvVNqL0D0SUw3VYHOd7Bb1FIua+m653hJgv9ssztFAO9z9iII8RDCR/HmlKMOIuVWU+lpwV
g0otOEXzcyrusvfEYAZZrWTIHfzzu/omgdetFWRTKFpU+gCh7ASYKtMNjRyKJK3AEzuLi9h3x1/X
o/trFY0PtaDtsfiOtY/CuoJoJX0hZBawehM2mNUxo4PdWHB2JEZTm+pnR5xqqZE1fwzgBlw9zp8v
H8V63SePU4zJlu9dkCbdGrc8g+DTJTM6AWVN4RYsi0+7iyA5Z0MTm6+59deyno7Tyus8zWkDsGoP
X1RchsG0iGuarGgFkiDzpSBl1GSnOQ0PJVaunWLJLkxjKO8DFkfazwiG+DnWu2pRXefDilcmuPut
OkNI6V1GSs6DyLrp7LFVg32iFd0KW0XlNy/QIdDm1H0cR+ks0gsTpW2OodYGb6ljANBtYl2bUXyu
ufIA7ozFNJrTr1aijlHOJ17KuvcbvTMyLds4LDid/ssTJpYvZZoF9kcv4qeBIBseXiNu/vJDD2Y7
a668xAJ2aCsGCe4A8IGFaxgfpifvu7fTAdMHbGsLq21br8FUJP1Lt57+9Oe+FcwtGcaIclvOhltm
O4s2V5GlkaVamms1DNUgd9Vbd5Xv0EGanxarJSmHeFWyYWeB8ojwOmHvV+UskJhkuK4fleMRlvT0
VFbr106nghPGjNVC8OGdjOt2RwzMUUCavv3JHXNZJg38Em5FCcYlWXlbnyyXHMkLWJFGpcmFYLeD
mIElzP5ZwCRr+NXHH8T0AI0S2ZQVv3e5QS6t2FVFVQrII3DFW5jYVYIHsx7BYrz+Rv0vOF/ZOtw+
9gsh5ARamyq0PKzhrZXJU+9ZZrFdRtTNQdaIqNtTt4Wpj8I99FKmj+9xaniFjCE63MbPf8x9tey3
UAg2twOrwzblxawhWzn5ZwRy+8Ig+v/KG6Oe2p3Qv/7hYSPxX9DjIwXudEglRQIKUKG3kcEaZjmJ
STXw1F3PzXO0n/W2a43xJjTWQNCOlt8PMaPhW2yEhgdDPBGeF/B30x+oAKSwwYwsBc0HpB2q3xo7
PQZuYlH6jODwBu7iL/bCWaaBSQVzFBmTyAoeoETjCwB1SZWsI3gIecgqaCfpSNwpkm/ZqPbXHZib
5IwwoSRPqS3qyk6Z1wvPkojj5lkDium/yoVIH80dvNcXSSj0Ptjh/k3W+JxkJWEw3QNgIRPLnuVV
jW8XNA3uNbOg5emiMoArxJymAwBaWHDCUqCsQlk/DfDUviau+DjFYjLyeI0ZzWpoTNg+pn6CD0lx
0tX82STNGX6ePHQfwAkHK3kW9pW/emGyP8ShyfffQTl712JK5KqgN2xgmgsVACbA2nSSFX+CkciS
l/frQ4lJRUctlM0WzxKtSBDXKkf628wFa0FdQUAKw0k9W3oW7m6QGNQeNNyBmTtB/pr83n4YmxjJ
c+K1QfI6yDIyHGOm32Xd4D/M7818imsbzpPQBlGEBdaVgq79TV0vDmZcjEvxDK5IuO6NVM/2WB7n
+51n+OwKH0D2qCyHVwnK4qBxBM5cobDJnnLvkvqPGwWrkl0Vw72e4t5ESNSnGhr9MXEhqsMz2TBp
hxYH8yz90ABZ+TdBItDyCY3dLEnlqNd0zGCfI3jm3or5qX2RNjp/bBUCYBX4sSpHaDXNIGWxurZu
6EUohPDsOCIBnyTn4qqGx7yZfMOxGOtQD6srQ9qNhOt6GQJOmbZzyiF1c7DnFgRSTc1bScCBBv+v
uPcasmPUaSxagIoqyaY6HuvR/QILb+0O8hhJiYXod0gUUGB5t0OSK3WA6Qg31gJ/hgHk6PWn1uhq
6UjnIuf7avKEZCvU6NSPGRmDKnzly7pIuowQPrbxY4SWT0Y+nglEpkSU+35y5U9EjUPF9fQq2lf0
wGLvAJb5jKbkPik9DYWoMW0K0xHSlimp9bvBzKXiPjFXVDpcaUqOvPTNevDL/3ZhwRsRbjedm7pj
OalzN1IiOp5F2fwj2IhFIEVfQS2m6kUJXUOBHXIeRgaplaKFb55rp6y+qmQYWSo/HOa5LzGGJIwb
ZcWmKDIfVhUA9Qu9D7j7Z/virQNu2TvIY2H9pBYORhiBXDr0UHeSNyCKnNCe3sfiXCANtl9OSazV
bvyeQjbDEDnDZUp4fsKgeHAKuRsHQZwMVpE1Vkxln0Hi9MUYJDTHNQr+D2mYnj5CbgvKEUdTsN16
MRMsB7Uhk//5yHaE9x9Nafh1MHlHTPKFG0PxjuPFAJRwROcYdFWNanZTPjUOWZz0SZ7IyrwMzxLt
TZ6aLF9SaZohY5qM/ybVstLLUWnG/9aFPOSNUVQ5bCWH0AaofLeyh6YeqFokP/8gVskPuFCz9VMk
pvl56kut5yTVj1JDSoZGrreRV/XuiMSTcXdiRrmXUmxAyNkufsKXQlgyJ9EGa9j0DV1pZ5yckPyK
fj7XoHCMlbRXjs00fJ+d2a92NbX5D6H3dKXDTSmT2avRdphNeM29+PWkXsYuiK0WoBpjsIX4mTDq
udiVMW0fSey03uXhn1AKEwaYoyC5AhDtVtL4ckC/k82NrTw9iEVvUCUhF4VwuhnbbdJ3o31Q9Cnm
od+idI6pd2qGLEexfn8wJf6KdIBEdEqJO1DL8gYNQvMHigX5jAHgzKrsApbKa1RL8ea/OxqQxspZ
QBAoLVlkddWQdvtaR/UIzWNWYMbEmF+/bFDSiyoICjBUIInrl8DJ78EDIL+2GA6nEUGl3r/9Ops9
O37chWVZN9BRnIeYpN6lJtGlXdhejw25oqrahPAKNdGyiV+HV5Yl2lnLuhjfmolRqbotpoNT/mJ9
U6qRGNpOtxl6MvpszkGGk7wKcaX3hkIDdyiSIYbUxmDXqflzZVqjdoRYCvipc2T0WKb1L1Vmj4hv
9E5Gbp7KUrh9grmDpbpcBchjYBQqJ5qGeOYJQGKh8ZL83PHwB+zMTrJgQLnhqDOSHtFd0yx+CXgk
4qTBVDEmRnJ/6WcGJR3OpvUJM1O2N/rSAlMyqC6zoMky3LyXa92Rx8TDIPVgKnh6dvS2PiiIQ3Q5
8iE9yBQ6EjbQAhQADb1n+rNdCduut/VsrN8OPKLwJRUkxnnuwli8H+mEAegqHeDXsqyVFvUW2EeR
OtOZxEnJmN17WlMprwXH5PCCaRlzd7V3VDMrb0xhmEE11kWa5h3KBDmk8ISPlUXO22oKPY72sZGy
kzBTVEFnj0moqfQUMEY26G+0M/aJBT3gKaVQsmUBGbqYYOaL2RB8RhjSowgKETpk3e5pT4h6NBH2
Lw7E1oh+XEkYCOnh64NzotN/k7FPg3EZqRMSHVfj3TDSS+/emgzOw+0WW46vCri7HPC2v4YAsZ7a
8ICSo8zxDkvPgrUm96WFGqspimSz//Xf239vu5Z4gHLEiB/qtOM3/kjGqou38wwxp+UWmKi7RdjU
PensZjzPnfD9fQoKVJoFSR6mnPoxuPchvfUWqGDjkQTwIj66DlFxXkGOybM6Ht06p9EeF69X7jCm
kku9Y12bkPEznJEETOULF0o/HmT4v2AkNcndWmx63UcewG7CocV2TQRkeWiZ6cXT/T0ROPp/HJu6
XvNm1BfWcblrs9e5JecYVV7H4nDpU1nn6+XL/eivM2rAyzp81EOZDCYtrT6ONoYPFq8eTTR0EBoe
LcgjjYu7+InlgVmB5NkVpjYh7UIy7C5qSKl8vvZibpHt2iMfq8fbW4gRMOJfNmIJi3cww9qjNnnr
5cXVchuKGNrlWwd3xDOOug9HdDeZ9UDOMqb3TcQjUnFVOl5O65O7y9hx6ihwo5CM5ZnO8CO2eNqw
6GwiuYPDEjDVbe+X5uTESoosfwavTOdYtvI4HGFPG5sZPCv3hD20zBiqT4qZbQZ53zLEAlUCq5GO
66A/Qa6XKcN9UFl8WgqFLJ+L1i3+3Sa8nT9BebL9olXAnCGeg6Apd1Y6dMMz45T/m3IMkHJxOiF7
lzL+w4KFvkslJBGMAgcP7pJ5lrvlMQnb3fS8F7Q/3pN4AgQbfRnSwVFNNOYYhIyH8TImyyAnn0fj
/B9m1tIx4Tobi9hyw5EMsNGzPMezf2RxeWk/+5IfiEsivUFzxCgg31usnH4QDFIOsRUE1pfcfw9l
7uZIcB5IfPHrv1AYGb/+IUUxkSzEs5CIeBjQXjsxXQCqJlaMlk5zfdF0idco2MZmnYrr385ABtbr
agTC9WAfdPn9X1lOWvCgkVW6+fKZP1gb5PHomsIVj2cMbUN7Wx44qHzK4vRszmi0Oaww0NFFGp0B
tdraNVMKvXd81gbPc1bazqs2fpzqKuMkZI+2SC8QObjsHHPNTMfGnSh5lDb3EgOxPrqAqmCq4TXP
/RbAaxOu4Hbb8W4bXHm6WVyw5Ynn1ObSg0tEXaevPYu57Co7fg310haRGUd483422NpVMyWiq8dm
rHY9DFyVypu1mGPU31uX9go0VLOMHEKFmajJZDQe22bFRByagxf5AoGZh0vlApGwovkj7KUX5xR0
cV1mTAi9BJuWz0XTYJpBFh8CIBKnX2o/DNrYpOrs57CLonHhL4/Z8aytXdt03EhyrYfVhHYZftSG
42hv5GvLlTOKT8al+BF77YY34XRaqiYpaSB69yIA2kR6JjyX0aeu4kIuXMbyMtxbCQQG26yLtmlx
ApkgHiNMoWsglmghT3/A4WmrXLKEk6FM8+2wbLJZn1Lcb+0Axo2YyUDQdxz/k4CeSHSW4FNjphNa
pPeD7yAR6n4FkU90MBSQk1DjQqNIffHOdaAK4z4ohxoo28gtYLuS5gLTH39YKbR+AvX1/Jger2yw
78y4+a3duawhULdRpJwBM20cY0HdNa/W5jygnEiY7caDISTg5siLu7RamkpXM6tX9BLMXOURX/IA
H12yELIbIMYvOqPgZte9juyBilMeaevCXZj5JH1yHTRyzcTAvfqAwGpMbobTMwU2xSgJ4kbRUUud
3/a5a6hixv83OGRAFk4LG59BSk4eWkt9fvSTY2RJ3b4RUEzvLIzWYroVnah0EjB+687QBaBIoDr2
p9LUS21jCBZUrUKgrMoW8xhVPfL4pjI2x8Ch7tihPchOFG+talIeLF3iAKWjT04EtSFNsOYR5NHI
TBuZ0uySm6hYwlitEBZsNbTSPaz8kEqFe0LxaSL2Z3Iy5+5JQFXzEO1T9mQW9haKztl1ZYiHXMoc
5KsS91RUwwKuzE5UQt1EfbMS+iQvnm+/S26m/wrxvMnpIDb4iSwzRHzXbw3dg3kYwn1BaUP5kCRB
q7AEH5p5QL9DsNnj3vHhgmWQWo/K+hfBQCuiFj568+NBG7syGvpXNHaCcNrn7GCueP06Dqsajsjq
o8IqevniCgQJMybJqll17kzVfOBLBigL7XSTgDKlr/jSoGMlLfJGhy5Okele0xWE8RjQsKXtjX35
iWY3PfxFzT6ZjO0YB8sX8WplXeDdygadvIs+CAyS8IEok5VAzYQGyUvlb42Wro3vQfai0kohZrlE
shCGbXrrLPuHV3o1P3+WDND6A78yjgULhVHVDuUnudgdKUh8e0kbFLYHjn7oNKzeQ2p79AmxwI9I
yZaUFCUD1vd8bY6ErZkOnHR0Wqy6Ftk5K7IJpLrsg8rNRz9NLz/nQGG9KFS76ebDT+NVxq5L5mnm
cVLkwtUmFVsWCcNFLVncdJlz9P8SM1qdnaLbX8di2r5JSrJWJmzC7MBXYa5sPycaN+lSnrxo0l8N
dPhwoyp/kyit0aScCfaZkvmJ1gtOABJj5kzmkk0+IzDzhnYYL15YRynZq/pMGBqPct2FKdvx9NnC
rkmo2WIWRQTQ10Vsp2ZZX9CnT/0WnMTvvWGjLb+BowRIv2LSXLutjwpyBPnn8PuwNhomT5/cjeRF
YC6KW1ptfOUSmUToHjrMeRgztFQLZQzDXtaPpY60V0LHovSgx3dZ+QLy6VQTR10bYWlATAiY+Oa2
NYkYYKLnyLrASwArRwhBtKWI8XSJ3TfsESJgiUkw7s4oNnYBlLBEA/LGLpZqWggxu+7pazx0FFnL
dYbcFf2Erp6NwmatpYzyY1RS4/1Yzci+7LkXX6ytteVEBZBcY6JTRM1srQaxF6L6PUN3HBtzh4z5
OImBN4LTf6H7iLwGksUZBhXud2ZavfoW025jbgQQJAHp84jVkUTbfUidws6CA5VxYIJW1E4Exa5o
OBaD5DB4bXM5kaVq/tVfu5hJcnDioLl/H5p2NgXG6ePBlzBE6VGrJD5KN+bhCjUjwmFe7k5mfIlj
pasiQzTFIvmuhIpWb/veeSme+j8pSvWaFwZaYxv9SLsgklFYfd74lPalOu6jkwiOwnjXSjpO8d69
ghjr5H/CEh4wn2ew7WCDFT579Vc136efWSEPvNq796l722lB/RrUuej6YGmj7u8t35STobzd+H01
vdnhJAPgLCMi05+ioSWXqXIjNTXPNbsHCvFSldUof8K24FjeSMHrthKlheqZsPNKweCezaNIpLP1
7043MC3/Zif7NKGWOgLVI36BamlgNTn5FzWd2uA1vPMn0SkZPo6mjaXoF/Kamoe/cKb/hllop4v3
24uYs39QLTQF663jJE7VtZ1QarGyW4bU5BL7b0VB2/x2YjPtIrH6GiJXeve+rbHXFNEopxyZcfCv
jxduJ4wzmHWuLdzh4mipwxXCzy1zg8OCrcV7PASiFw3wswfxxfjs2Ud2nhO02EIwgIq5XZTet89+
Gfyf5UsQl/mbi32cJV6FUI7afcDkexNYTBDkrD5BX+4vP7Ug6X7hY1ZnkO51aV28GQRLd++SP8kz
QbiYiidOkb0Kp/jsrWL5Wy6zf8imWOhcZ5LP7dVgfxziSKa+Tzi9XxymCCzjXdbTSKU9sMhqm4JS
1vxbZb66v6LMJZbgFVaEAbFlMP1sXbaZsmQYm3iKJF5/4MrvuHHEnaiDg7X7jlwyGhDYXq/nzSRt
jSxck3TTYP4Cr7+DkIDI60hb717jGmQ4BP+75O9xrmprQ7KWl/KkH5ddWLMlvF2BgkspFybhvsx2
U5Du80PXtrySI+6eeYfpKg9TNYEVBZhz9+cI7dxDCT8kQaa6hgxTFj/4HhaMHQyZqQEPQJ7D+AX9
JQs6ByOyoh4Cev9bXJZ9rQ6qEbQ72OTDfYCXa44Wp5Z0j9BGn+eTkDsqL1mUGfCWPGbDOyZKaunO
36WsW+5A5z7lrPYSHU7Kt+fr2l+uhB/R3tK7/yKhRP7LPufDm90DVCDKBhr6qqxxNO6+cqQv2him
TIek3hUpcIda/4cGC5PLkFdkKsANLi+Ea+08qkArlegzNbjnziDlOCfFFMTIBta6I0mePwAW/+Pq
Vp3crCGrbwc/d1+sajkQccvTQWMxwt+KGyUDrXcDVRZubBvQkQ8sChN37DIgO8rkA2gHTPIsCq6z
tWprHmbh3NbJPKpx0oO4WQSbKWR8fdmU3yPRjAl7aMteo27j4yze8A9hxnMLRub3GGvipBHdUQAk
eJBofMRTTJg0QMxshOybIv9XssD0+dlWKKsaUL/Kmhbj23a0YRWxQY/fHuLgstKy45hEf5uLlCbi
Mi4ZtSN4VmBbg3Q+f4huC4FJJ3Dc+3l0ijX5HRqhS7msefxzveCgjZ32XBO9Yo2FAE4m7oi/FntA
oE9CwaP/vBYgs2ITnHiatj+0Khuxasane8Tp6f226zdLwuG0DP849DP4pis4ps23Y3teVBiRzCjL
+zU/7MmbOzev2441iXn9lcD3NyDwuuaYSliWlW7902HSTGCpls6XSwdxiNPD4hPJGZFabs5pwHfF
x1xzDiE9PNGLjqCLN1PC5uIBH9U+qKuQ8q/IPrGCImulqeOiUZ8x6R9jmqEhB+NZ/dtQcTo6cczP
Fg+eQCnd7wW4R2uCh89tqtABOhLtyHLjpdCxBBH4KAlTjH3KT8wdVCQ+Uvva0Xs1I6T0CU0467Me
OIGuqY/qiWnRcw1Tr+QfpBaxObCuNN3A0+vPhiwEH48CP2liHr/Sia2CzM60qxdXoLUT3RhhIgjy
8t1GE9Mbr2lwcuzwkhHmXBOrtW+wJe6Tfr5IUlalx/w9ZnkfqYrPIvxiK/ETkf/r0ajTgOCxbpWH
YBLiI7fuaxKpO2eRDno4YIS74UktN/9bLVEyTM36TdmyDoZHRA9CtVUDJlpxDaTP4EBam6Si4AyR
bjpiug7Sd0zzBMjsBLe1rFuT6edftXf7297z6LsJLH/U7HcEcsiNGmbTuBcgsf71c+SuEN1pK0rp
UxM2dbkHWwg2AF6ksc1Hek79aFT3GzyAQNsKLBsg+/IPsyuRg/4QlO+Civ+ihOif41dJpu1oMQBq
vl08ydGOpFJl39ETNSiKCCexEUfE2di2HMIeoTUMz2g5xnpslmxsBj1OB5LawrSF50hcCdEqOfnO
cyUhuW+X+gTgEhFVi5qEJ5bG3khgI2sik6NfMBwnQtQHksJ25LNrJb5jPmDSaEMOrStrgyyj6Uth
bWWnDmQDCmjK4TnzoxzBBbyOWnNgQePSsZJ2Dl4/qSHQpuecxR0O5jCgSjv0GBOF081CTIcBRUZw
pdJo8PlZMtBnGGUFQS2Wzt70JnGsWIYgLspWBImEAn18Ruxi/PULvtv/Kk/kgKOUZzBHrCL2OQv3
5pcL6jLpjqRwLY+JBryaGCHQnR2b36YFcrPZgzWmjQNjosMB7V/mPHMXJf8cK+vlxA2kWyYFyUGA
lkV1DqxR9ni2cuh6+uKn8kbk4HzB/Q/cpONEDiMucwOi+6YiJ4XBm03LNnPwziSj6zrOPbNiTlXj
+mwguza0EkBIWoLR+yl6p6zxE3GKLvJ1xiQscJ8xiJuiJoEr0vGabKqYA+DfZTLE0M+YIUs8Jy/P
rWx9F+EGIL1kP+jWO8JBQe1+2SlDI5B/Yn8QH6hxW3x8TdDgYTnEJ4oWt2tJqhV3BGMhI3jA8e9U
o78x3wUKp8GRUnub/nngMKPRG4qMX2W4BNozYZ+8DdUMoQKhgdD++dBiFXdGNK40g2zIfjJgJ4Q0
uUiJtkGac1ELfOPVC88uTjV4D3+t1KxrGv0bRkMcRwbqyrWILMt3mzbB7zacGy5ocA7Wo+PQlSM7
GxFs4vYh+96a6qai2R3PPEGfu7+yKZHhU57pcJd7Q2GXVS0pXOWFIOQVknX2ocWl1PGAlRmDBXgX
8nv+P6lLmT0zMynBO22NrpDyzl6NKndZPd3z8rGKy3TGRhVJJcfGw5+jzqyqbuTFdxHbLHEnJSFT
g5n4aIYBOhYKYFQBMUkWHDGRy0dB87XUM+E9rbPZpZ7I/Ib5mCBmNQHogptU6W05kaeK+YIRolMx
SJKAWbphFae00Ef3ptYW8pZrgyBq6vwHdA/exI5/bjjsaNcarMyuM8Ql1g0o7nPd7Q9YbPT4ovaw
XhMWShfYNV3oUMiwXrigJmqzul8L8xyfC1wbvl/cQByL63hV13TCu7+Jm3jm15cXCfv67a+4HwmP
VSPVjL/ezW5jn4GnPCfOK/1LyRvkc4vJj9Ineh4Z8vDNrAJe9DUx2jzAQClJZNlt4COD5H9DO8f+
2M/gnrU1WqEorLDpBzcYEXgJmRase5e/wonDf7jV1ErKYrBbFWH0/z9IMNGZ5xEkfxlTVXr3RnsC
7AbF55kMoZSuy1ouvrsZbJMinKFwTyAUgm6frEsHxK6j4+nJ5RZBwiO7jpoS/ZNqhr77FlhyfCLV
6M6ZPsMqoASkwqYnjRZ/IrFYxDqT1H0VblC8E1YlnlXBqk+yCcTtJJKQM5PfqKoz0Hoq6C3pP2Pn
Pb+1IStrMUl0xmthcKdGm+3C81jUrsPvgKMHQAta3VLvIsAabSNq7WE26l2Kg4vRmN4d0RvAVW5J
4hURFnzLkveQ1wJbpxBOylNdc7N5+kivx789dCa9mdS+y5ZQ6ytexx1nAGXNdumDJ86d42GVIRGI
5vaniLjRcJd0qT6KWUNIgd+R2BjIvSIkfXkByz4rSeyQ3DWgfMtRMAetLEc1W3G1nYYFQ9qjb9YZ
3VfJmu1j+Cm73PtFIZ2nGb12LYlB9L+2vki7LL1x+7DnK6LZDrhJbseeWFzqegskGgUHDZTX7/j2
bHr56LkSs1AiX0qQC71rlz+wWoauEts6SVtELEjBUQaglboALF1zxSl29Ahk9iDu/wmgWzThuR9b
igbHObHXdpuLrU8u81qTZvJLzl71429uiCoT3pssCKjgD4fErVF5carF1ZXvN40NFHKlpeCBkdmj
PMVArT9eWGAzUkxQ86YUXf7qDbyfhjeYCGu6BmL/KCJJm0vXN81JbzdNMVbwRvhiIrRgOeVYAqst
kEWw6HiwKTRgQX18OlLBtQFPBrpumKNFsHIWbcDSWbywgsUrc6Ix39rMQPe1reE69hdJbXOKgEZk
1FiVC7Q0N9Up9j1aKiQO/jUpW8TaVYa6BFYAHpC/6S186ooObONoWtLLFdNkvq9bL7veY7KLlTxe
7I4uRvXi41Gf1XpWeZ3WNPP6n6mjEXo+nf9SEUuXfEezGDwwtjAH3RoVyy1zS8Uq6Tb8rMALC66r
JMoNVMuGIp/xRcDKCjGLtBabgZo51eooNb5ngFm4/xBcty7uZOqB3wmlneLkj78B6jL9NYTdthbC
GYdCLKxsaFdp8rwX3UvSJ+fFwJkzm6WUZZ3879OJsIJKSV1tEvOte81wm4K5GfUQRLz5a8vPEu5p
i9LcpR6H/lqc8skSgY0330wAwwEk9jw9/av8jYGGlaPZCVkSQ+i34HArFh9AgLwFSki0+b9jjFsy
7MndyQE1bQphmkOA/FPPsOlzMwiOb1V2nhsVT8FGHu/p+nAcOwfiFKGaLTO0wLZ1nACqMME1I0v5
jQD4Np0cNjn/IrGxNaYL8azO9jCN4NzDgnOm5bBpLYAlxjSWsW2MbRoaaaaOXKyl81Hw8gC3Zw5h
x1gvm+PhdDdfzHFat4CPUvDEgDqdnMTV0XyT0sd7GgOqTqtUfb3s8c53iSdoJ9P+SndIJ3Y8kiIm
oRfcJ4jVlQzjszccg0jL+3r1YsoBpX94InhtFAn0pr+eULAAkfOcMrhXb1+8Cu+Q2TkcaUx/nsI0
VoqMZTOJ+iYCpv/8ZSZVFnm7YTqjPWOlShWRU6rq6NewfbAxuymg2YOjPG/1P78+Cne9qbqELNnD
GFMycQnPsYl79FSU6C2La6MRmlf1bmsWCdFdbdpD92kMkyFztLpK4XyQgiWEPWbLKZ+W1MnuaQs3
f9Zb35A5D6OpAM/TJufnNQQfjk9wqIrwZXo8Y4bQ1wduy6HF/Hcs9EariVPAkial+ZqnqvjQEWQ7
KdTmV84QN56boyRjnICPfvwsjj8lApGgJfSJ/kwlyxBBRk+OgomZpQVY2Lm2TWmImKqJlrVLlH0p
TkIBdTpPE6mEt2kQOxBxTor9oPPm0rPjgbOVuFHYTz9MQnLhiTp3zbcE8fBQU6kd8fk6kU0Ve/Qp
90x4k6YCD7ZAK2auM7LHhdV3l/H4wTPxl0UZR5sAhFiaqUYKs2mcNNK35U4Ng7YtGjYX9179dpCA
XqZityt2ozGXj9K2sbs3qqVbfZ+xx3zSRIyQfkIPRSTcd1b82NvF+a9VPL2mF7aiHQU+7rwUtmWI
zxIqyD82jWaDmIcw+gR6hzrqmiVUSeBGfdtEJnwVv+mRXniQzDaJcTVj2x8EwutvYqQsFHiolvxr
2a9Oa+AXTkEKgNs1J+CGEGhVP69HZC51Rcae91sZRDkjTDTfrfhCEHuFkI3eo/2B/4yygTnW93fG
V+XJQgClaGXDdokNVxNtzhWDw/1ReE2cnV+CICa4g2CF2hs8wTb7nnS3vvOIvU16M4acGeZ4hvLc
njeUwl2sBD7raYAI5Vh2LketEcGIMpbDLWTyJFVKVDb3jk5GEQjTXWYn9CMcAtASHZ8DWDKxWx+3
Fk/UJC6ck5N5DbdehKyXKcC8bNcWbdSvpcLmMvviQgU9g8C4Uuzssv+8UVnZ7wCqA4Aa2V16ganp
mgbWDtekOwMmHNiIvhhdAXjUT5PIrFXF0UaiYPCKJTuDYgV5JlHthd/LsF8snNjGCrAIatxOslsu
PiFt1BH6nkJf9/abfABlonEMlnj6ex5wlaEpExLRpEgdQKoqrneusGl3j2kfKA5IjWtxk7AVpQqT
tXBHquj0bx1Bph7EzQXoif8ClJRAgA55aIMATbzVI/uurniNi6B0ChSVkmU/YOnrllTB+cUk8tbc
aPHFwyLwu2iQov4q0KaBdJbXWIYWrSdRVwv0dQqvvWSQMCoHurkpZhiLlawVF5A7/9R+QheQZFU6
tCtnOURZOky0gEZfAPoIdN946dZ6m4BQOJdjSwrqBTAqW/Ahh0JkP0fNlzg05WroaUPBnn8C0pZR
faAKW3gOx9CJwd8b0Qp82hwm976JjY+C/IeVa/rBH78Yl9GFif0As5ekxYxNkuJk0CLZaQDIXApN
+AWJzrXUdoEpSbnUGUL8eGYbyJ0+F0N65eRQytgOR1a1Imy4HX3oF1hl8jc0uqR5NSRzcZg1EJuh
jdLWDN8NQIfsuGfhE49MxI58RD58UxRncEOhWcHeheJewXalleYNEYoFu2sieEFx5xO1kJCUUP/8
3Uc+A+UjCzQ+avoljv8GWCrdSejd1wM117nRV2p69nyYo8WxkptzSSZd9lvP2aywMs+nK8HilNtd
y9d3pYgStq/t95nsR6Il3OuGzstwAsaOVWtHk6D9bKPlCtPA6vUDZQvFZ6By/o/j7qorL9PhtpJ5
H9qQcD/mZQLeCCmCF4TsrFQ/2m3bjnBT5iJjnhdwHxGulffd/ZalqYb3zg8faMtHQ+hHeZ/j9w5y
p17noIG/+tQucmgX5C05SiAYmlLaoGJIB2JjBkyPGJrTIma8DbZhwk/a57P31ms+Qa6WLISjCJUd
NjHPx41eizsndbyGc/F+w3edp0MySmnI0lfyXWZPzq4EVltvugKrDicPvNK3IO29B955SzBYJ/Dj
4F0QVN4pMgxa4T9B8fJmC10EmnviWfwCtgoYjH2xIiCNEcYgOJlDQC1Vtt8Kqo+q4ZtuhWLwe/8f
/wYq6gphsWaNxe9c5HR37FOAfriP4ai9KMzdrj+zKOSg66xDB0+lXiB6xtu8J04pbfMx6OrBBuYs
Apl43ixHZcTpfT8UGpAW3+JS7xhSoUjeL7CwZ/Y9Q+OacsMO78Do6lLfkoPDGoSTfQtlWlx7JETd
B3jFkLsK2gsQgKo8yMfgKQNn1dmCYtIbQPncWXmAORPgbiOFXM/I430uGOOizYkg8pEdGD6KdJep
CbKhXfdfEePmk94JAQVpocXYvI2xsrt0/tRRpC6GfKLT2vuklYOj7A8xCgtLFzUUVsFTvoVJIyNu
BPbQk3sMPCIcJpD5QBo9DAQ7Ko/+D3Q8PSv2FN8EmgQKf8GN+AtD264ShC4lxaW4jeugyqEJjem1
3t7s82Smh0zBYwBsBqSLgDq9lmCVtZSbyw33DGfhf4CfvSiX6GUbK+s+eEmhw8bJs1nAce0qaotr
4uT9hjvBfiT9CLVyWZaAUK/8CogQ83RovgBPwrJ++YJGH8hGhyZEGBbkDiflhRSm250Ot7Vy0v/f
rvkRtz32N93X0R/uZEiG7uuZ1lK115sHv8+6Wzx+hpkCJe+vpOqoiR2rbHm++Q1y+rbufqn/4/WB
fImuuGu2v3/sAO2xiRpHXEQNWeCYBQdIx5mx2K700trUcennG4mqHl96Z02pUW4mv0Zdr+nu7sEh
MqsOpYOypA5mJPI70gm37+//mzsPAmuUNNnNtEZIYB6dJqbId8XkNtZMBqmi9F9kUk+mdGCX3xzo
7C1CLCyI8qTx4Gf/5IUOxpmUbjX8GqMqpEbuSiJhUtpSMlwkygoUwfPDoaSmjXnCBQRXahSzPPla
QSFNVKRstaIUh42awL7Ua3MSQ49KYmMbjP1Jki9K06u30d6Xo1fI6f8nFcT22jrgGkbVwRhK2uw/
ILrtaU8BUIoiM/YWVg+hYJYgp2PB3T29GmMNlDVOhxMfd4APFW/v5cDPN2rqORFGcLE18HpDsVbZ
EN/+HzBYGl23FKU7w3+6M/chNaFtwD01J5GJIsVgEs3r/4ti/gc0QPH1QtOrv6Sml4LsXBC7171O
kPchEW5EDDMan/tV1ZrLV44qoc8qvLco/KFQzaUaWm7pIMHjlxI4HHogwP05PuvHM2XX0kLw/6Kn
QTeiF1A8r1i4kGnLN2TgQ0wweN+NYtxdwjdQgsU6MAMO1qCRZKBI9kY2csVg+EBXSdK7OttmF/1L
lKOFg++eCy4Dr3VAmxFa9/YV+5ByQSIJmff/HN+ebExooucISSLn1s5g0br/G/AiM30wq4ycG/SM
l16ULQdRGRDP20SjDDkcp5Ki061Bhazab85REvD2BpvWTQORY5r9TOGrwoPwkuIohGT5PR0yxC6O
W0uhNqs42iz/TPqI6QH4dkbY/kzC9DceQwQylsQyyE8US+vC64doRjWhF4Yi8H10Z16vTKu4/p9d
pM0En6OoAlPRaPiUo0K2IhHF2fAH9U5F0kChxq3EvMEfdz5XzM5SBVidWdZ+Z7w/ufNTY5jehwGK
jKatby0k/iIujLK/CwiKIga0DG4VT/Sjd5mJjZcEl1y50UkeOgX5J1lk0g6nKVh/D95YbiDTLU7R
o1MZgeX0NX+8mY1RISHLXIGupsBRncINi98oxGoF9ZOpDlKYCDHN8GAnvK4MMxeHyiNLoXbjYoA3
ug34SH6kpXWBA9zFGsyBeanuUlgXaBCOvi1JDwCjy6/kPICdyadCYCbrIC5f4HEwSe8LVyaPEpF/
FuD6MeC4odkzZ1+NgSMZn02H98+h8qtBHQvpvoe9YBivMimAJ3R9VNrvnMXWI5wSBuDIQSEXZw+c
Uco5z+tzaGc4sw52BJaxrsWAarjJ85cB39utmMwMqLjjBiyGxE/LGycSDNN51CexAkouRrQPQFWg
FkmrMwclveiETUapqHpBDE4ptuQL6+3Rio7gVAp19UV0CVqyLwQ0BjjyXV/9FsWZqFwtUJYsKxTU
KxS0L1hipGQJm56DND1ZFW7dk6d/wDnEw1IRqGumwtaZpHJ/LssPLJmAWIv0H/o8nUjcuQ5YNuB7
l3B7376digz643rda62gMoNeWMouiv28xjqy10ZeFjkbBEFDm1cy6zCD+epON5fEa3WkBHyE15Kt
5Q2gJIwMn/TRqBPUYkhGQMq/uwwDFKui7w0hvUNateEXqfQ9bQBhCkjbyFd3v5aqd9q9pj4T95u1
dw6q5qDuEe3fUXDuTfRt328XpDPypM2wwVn4cSUdrvqrGg4j2J94yUu8QDhP5e51RjdMLXinB1Nj
k3qq3m6ZHdjwchg5KfsNdOFtNHmA+iHIP0EMnT/gNRJ3i9EHcgXOx10WS6oK9hYTzckvGq8LB9S/
vwUy5PBBF5MT0W0a5QbSauGbosDsAsm9a+bV5v7IikoY5ICgdhiXZg42YhUWg/sn1Tu9783neM4O
SyrsHyxojr+AL7/3AbJ/uZWriShG3/wOtJjhXKQzasvS5ectTqaX1niL6dVMCXUMrLgyDn4fyZt1
ewsX7sNFkeQfTdleIuNNSwR8Enyij4k6p0oD9wU+GSRAOoSIcB2VjmfrscKAwyJ02Zr2dGPoMqM3
GkvPJpTDouFpJzW/AwdF4oMFu0t0Fcn6WEtD1/1gJm5yF+Jqn03GaT7M6ZAe72VmKxsc8na0wGRo
9djjelcysfUfzWIPmr8WGgnA6n0lbHw7LK7NezbvGm6QfW9nB6LdNSPFAt30SHWEoRyBvQa0By7o
J9NKSJW2XYUGATIzRVV7OBWMBOBTUdqhQcrRNUbcocUxziyaxb5qJEHTbvYZjifizHQwZuHngNms
04d+/B/ehL7ADdl1mew7cpD+1exQAS8bFux+A+rHX2xsXgH00pO2piy0C7T5+fQ2CCzBz9v7ZVFU
7H8lnZtM1EBA4+sVyWUPUN6tjycm0aKFrRyAgxZZM9D31+JlvXIGXmhGBcOq7oDpo5Fbcm3VKg6A
SM5ljjdgXICzs+XmaDTzpjqK6GIXzwJFsH27fpxedHcXinqHve5pLpDnjYcztnUSSbN7ZaT9VQzG
Ywu2QhjFIs7kS1mT+ZFPu+p4X77p0gHm4IJOp2LPDh2mYuaOcVbleazExpvsmBYMubafgnIcSkgQ
SX1GZV9Jwly5Hquq8DmhwxxG5RQFmlJ+TBhOjNyFVq0M58CzAVbEiAL4uAiNPLGxwzhx1hbHr7GP
EQiOF1ad3BUb6v0Cec7DhPWmi/JeROw+32Qsy6mHs6Q3RFvm9deQ5N2oGNNJk9KIVEZprm0/H9US
jW36135/4Gn7gSMRTMoIgQbd/LqQl8mscZANNHp4vngdqxJxP51QEpgCnM4+izni1yrQyoh+ngk9
lzMpbsnujFePvtf/VkyZ2v2hj+FIwQL+7O7rVXKbByA17U+h2nN0USJhWhuv1T0GpsEFIHrGIhXp
myEoIL6I4hHTxL+6EQXglvwajYMZrucI1z3EUhDKTy+ln5L5lpCU8IPKslfMfc20EWTJqa7ztiDc
qazbsUee4U5w9x45BiT1FuZmPmL+m5S+uIKU2iXScs1h2pMqZBuJEZ2fCNtVBJOqFs2X+xp1gnFy
WwABUfj05VKeGGexp+4T3WslKiibF2JZjcWkjAlSB/1ekQlgfjRNq6G1gQNwhrDrN7ncWjeWrocx
qCUx62bJRTSV0UXFYFrjAT7g0a4TDo3+fCWVRobuiu3JFlOoZn2IjIsETbxo/8MdIx5uAICsGxhi
Z77CaowoEIQ68L6qhMJq5gsTKKN+QglNGRDdbbCpfInAcwSSuHnmwN1wsZFO8eMXiHv9xSxAdxA8
Ht74yFy1zMap0t6FTtMeL7rJRKkA9OWSMjr3iAb+9V5SsTJB+bP3xBQVHwP94fyL8deV15yPhKaI
gUlnFKifHSj2ixvSrY2Q9M8yybCzKwxAZaPl3sAqoye6F1Y9pXrgLDenNCcnIHgvvnYpsGtabOYC
c2b5E7kb+WSxcx6RADvJOa0dUKNsKWQqoymE3Cq/fjpjwOR2a/0QqXcnxzLY3G2sqGsXwCBH1fAE
0G48ftw0Q2kifs/ICydi6sH51s4KbGJS7d6wuJG6Vq7RZ/SeF+iVyIxo3oJWwWJWpDOtED/1qAWW
DVTEaHCMIb2YPh+v6h+KL+TtnW0sZ9Jvd9L29jkxdWGUqEixHMoaaxFFrXZu8Sgi/hgBAfaI1bTQ
2hsot29aMjj1N1X8xfCctAoa03k4zmcgM8QXiLJX7qK4SyVb6Md9fU2l5Vgr0W9HIjifdVZZwbOz
Gd37T35WaMGXX7K3bWQ02KLVF0Y/owCItgAdrQCIMD9Zlt5p/6JUgAj/u7gjtHeJ+f7D2Jdfvfke
olA4bbRghGMKooW5l5s6OGo0L2+mCpPkrz/bp708t1E/TtjHQjBU45LwDrrALGf+bQf8Qruug1kz
f/2ZUUJYMEeBVlRICkpq7W5no8pHjINxCC4NcSg1ArzRxfdJJKgrVf7+8svqgsdZkugBOqxq1G6/
hjSWk8nGM44fMbrxsKFZ7B2dxiAczwjtF3RcBKYLqF74ooCz+9C5WnorqOl2OGWwjiJW1PPlhvWF
qVKniAQRjUgK+FaLD2buosu8qPxmHZ8iRYlXCDgiPQIFZX03JTjsmYID961vYg6gHQU+oyHdr+l4
ctBzuQdwloA+hXWsDvHEJjzgR3C9NFOJns36YVx3qtTPJrhjoUgW7Hrr06irBFfvhcuATZFVW0xN
+CRLq8U0zrhoRGGkohF2VwtkKJALQRYc1YryIpfsmUCAEXvzJ5B+Rhk4xCRJZ0hf2tgH6BpoR9pJ
eSDaSo2xA3oMC4V6wYbPzINd7dBRqoTVR31DYfupZPpWCT+XRWF3uf90KZhOhn1TQ4/l5xqRBbNj
NnKfNa9YSCtkoXhNdSV20E1lmlQhJFBcvcIU8+Ts5uVm/jK/h7pWI1av2k1sr9pfa6fmv7zquEZB
qMiphVvjETHeGvHg9rQcdxv7b2A/hX3I1ye+A6aAX4/nZfbP8nbfVYauBu0oaUln/UkWXlBtziHs
9/sSB84klFTfPJ/Mhv+xTAKyg6HOF0AzjetUWxt1NE0U0K8ub3rY12gH2sia5NMMX0H5LBEz81QZ
cPZYpXC20MQ/cIu7sVVEz7cwUbp5M0qz8xhf7Rgcu446Y8O1iH3qphRXrfT0HU53a6Qba8MjuBk9
7WjOjfVbfk/0oS0ELDjes77GaJu46tqic0Uomn9T2GfPUbSFE0ycIELjBXIPHeCLvCWhFUTotbmn
INvKOfheBH2ugVr0abmoEHFV+QETUuGT0ihjOyTaluE0UrDWs4iexIEjJPRcy0ci3LeIWzxCjJdC
7cU2uEVdwZinBntAL5MvWAGZr9rVvQYmJ5MxiRQVSNoU+qz3TxgQiZl8Nh1p5VciiRrg6erkfm1R
G904MSTbWBh8fmBfgZjYcq+q/OJPD852ZJ+hA1S0RcfAm3JK5qJ+YCAlbTSBwyR+0doMxcZVkZeY
u3eQCVeY1Gyz1VslUzZxzH6Unqd1dkTkEI+0fqI74uHg9681vHj/VECAnWYDF1uLycWIAvTF1DWa
B4E/w8N51uLwD3P8d4ms34+lwd3CR+uxPBYw5k5MPhNG3zlnFJtU2DQRp9ZuzykZVIYlAsmJIfG7
HAjnfaxWugwQbnyTpbdd7dnB8NUqDsJmYdjiKwB4sP6EmSa//im/K0DNL2+XdD9z6Q8c8PTrSqMJ
bKi4ftr+eGtxVBaNOIVyWuOqJDASoTWlH6hEdoY5iMso4H1JPyHCVxdw8JEThZUR+Ufc6bJnUK2p
E83d46F13V/vektNiMBCaiHyj+2MsVgKk2qRwkk0h2Kt6Mt3aBptfnm4Keo2ncjFWIOLIaHnzp0U
2lJSV1l1vRx+uFhtpXwKfe+IjMXKz/pfzltHR/o4JUhb8FAaN1GCIeTCrtyME1Y+csRudO6v/dSA
Wikfsv3JTI5HsH/CM7Ym6g5qE0W0X5kHs8STKjTxQZ0QTQf/ppTbfoJlcnRPokixrBHG1C9zxsaZ
Jdmgb022XekHaT8LGMoKE0nJmhJZBUMRkNAfsaYZU4MtBXaK4fittpM20s8jHldS1JDMfD4YYdGc
Sk0EiRrtRLs7FEFLFgnxxNUWejP3WfETjBnnlfOVUWl3XuutYzjvZdigqSwh+1yrNyKu+5XfSbKg
NK/FdLtwiwdzeJ/lnkPbD/7JRUGloXnNKFt8GHeJZYiR6cvY3kP0XXJJSZX1ctNBY8OlfqVMFIBG
kzGpRhtu+0zoJoQzHzsjF+KCFWdtTazlwh6MvJSCc9ZB8ibt5ERKqs8LfS83PqSreoDGS/rdWxVK
R4TS8drgGN/0cPLyEfcpIMwbRoon0q2139FgPHxw9jYQrLYokMv/F1ighmIiSGG1Jr5oLd2o5nLb
Qwztwux7Ec/PHmpxNOgpJEvMuExxKIuO/Yl4Hjaf0Sp1k/GQD6dXHyyyjGZOcKQV1z3KUliXtqnt
L/KkaYAns4jD87FJFPjxAA4oZZBSGp9v3NcrT0VKeyk+R83lZhnFScgcdL8eBj6oCyDUcSLU7DJn
Y7e1YZFvr37MWDFMZj+jsKIsq3Q3Mp6Kxt2298tq0DlhBNwKfvZhE11lPMkNSpsk6DX+jFBwPkhx
iohYt62PN4dtZqePVdVxYJaiw6QweZRKkGnkMnBriRNd5id7KNdhKyQY1sv4NN+QCZa2L5UMrDNE
eZry8Sp+RJh+a0AjghFNOFHqGPoZZ8ZK80mk3lPJ6qCWIkJxeP98q2EwtaBSyth7RzXk8s9KOaB+
ZUIx2ugVkIvwPp0ObjBwwiHoyyZHQvcnjLq++walwtR9uPZ3xJOYige77jMUzmoXk0WER55Qt8B5
jwDg7ZtKpUXlKKq7h5nN+1PaBtE+4awkHxV2b6JOtSjNa+sa/4Nn1nV1eVxsuwvkeDc04kmKIC7c
p6Id75+wAUAw31wPb9AE99XSnFS8MuyiTNRjFE7ndg82KFBToYZsCLFKDkL7DY5QjcYb7TQNjlcy
vUFlKXSS3YSEWwMqwjChJ5FFkGY8upV97vdbMByqwVmCjJDw5FOHkLrVsA8rM+gQl4rjINtU0TtN
SgM4/0sjOBlqQ5zB7J6yex8Y+Iie8siU2LTiHeVdlr5nggS8rQOks2cXPjjHLSVtAL/z+GcDpWSE
aT/FxsK+1qEIkpOMK7JvHGEEmrkCFgld5i1oz/Sfc/ehiwB7LcKJXB2lxc/n8yC+YNQjZjjW9Dz8
oS9sSg9V/nWd/65JIfA2FtH2Krerg6Ccdg6h0PfeL7GAxazQY81124K5poPnPkllzJBp5WAtSd3Y
0eOs+kkulWyTk8jWwYUPEgODce1lcC6Dvpa5lmGAQUM6VXAj0bDTKwYrE+S/1wP3OK9WqtsbDEgr
UKlOBAuChSThA4RR3Klu5TjxJ42r9/DSwpe5Mkktg7HCaePqg+D741myy6RJZvelemXZQES1VKYV
nHn9E0xEcIpUERIx2i2HsljZOcME1KLDeNm9J6r8eYvECy0HYsLmk1MCBVZfq9dk2ZZxA0HkZR17
vN306/EVXNKWKNeL9h0VnK1enXXT5EjWuQR6oMfkbCtVyTRjwb9bNj2BLuLNFcbgGET3kEq2omfu
GfJGnzEXgvPE4cyWIKao8rNClV4OuSsknG8G6NLsENTVhGgkxS0h6KB3T19twJl+iLkMCARzSsSo
qEi036bM0NJpA4wbwZZnRHScN6TOenD4VGPe4fcaPNu4pp2d8vOOp1rsb8fN0Qc4qldhMgJ9S/uv
kBubyBhRX+HZ3RU2o8TXomxvToPUn4CsZBxdU3AjfSa8U9eJeP4JiSt+qKVtvkrL6VNWKoPhwmaV
CH4mDttK9N9Fxr1/Ybdlqf387Tx/5Q4C3yM5FiKTmCY+devEXAzMGt0JhFKtVweILD+7rFFDE3m+
wD3v4Zqc4FdM4JmbZ0Oxjkjr7WJKibEO4OixVElfbAUljuZNH0gLgD6w3rCA4BUAuWaeW7ZEO9jR
Gz33TwT2q4PDsYK6oi654u9Qb1QmnEtCThWMpml/xoB3rAg/x5zCVp6koNE1BRt+86PtPIP3HU8M
H1eH10aOU0pyFJTOiOeB7GaeVz3hFqdrTXkodL6jz42lAqjSIhVO5Yg/yf9jV/3YdTgA43RYCjvH
qzQZnlwLUJSh9FEUwFFLcM7miDXStLfFxDvx1oAxaeM4adtCxZ/Ilfi3ePy01zoZ43aARgXJCR2D
eJkagEFtHHoOuAZxtG1ASWYS4/4yU3RTxx5Xl/CtDT79VjSrdJ+GB7mzQR6r2VaVokTbW/kQJSa5
bUzpygTLGFNd15JVX9SZsY9iyTmseCmVer642n5ipZ/952PLKhtgYBrMmUprv4ZBt4Fy8dVpkBw1
v6I/oH09Az5bEV2zlNMSvmFBg+5uCqjEe/M1DbXJK7olFwocVS/cGvf33CsNBeYpK16/xZ/2y0jc
oEUBMldc2vDh1m/wYgXJCJu8mH81lRGKGC/vuyRj5iBh0Xbytk+z+qts3PVbcdC2OMI+SKmyXWMt
5ixhrEQUjMc7+n2GCMOLqLDgI589qjW9wjAWfkOSBw06UleM+ifqgoEyTOyn6HQykzGNevUxAE0s
mU/Fdftf2azXDsTp5fq2EHwniiWhQoGJUi83gSbsaHPPsWW87WnPEbM44QH3KVGTgff6IZXvPTrY
dPczLlWE4e1E3RsAuy4LVBU3d+3H4iPErL9sIyMLvRJoUPKAf6X1IGhp48XFnYcwHJzDDT1L62zq
xIM+ari27Dya5pjN8thvgjK/1do+N37kHUlTBuB7p/9WUn91AaRKo0ZhJht+yzAWWUym3kbzrLLQ
6izxDH4Fni3qiGkXvNjMg7WPnQjNBAtZwOiVmIZrPaMtvU2Skd3MZy5J4Mao6oW5j8caIIYK/K8k
hTL2xYk9gfmqj3roY9uZ1gTU2J+fv4HpNvtVK6z+o+tQ3X2zXg4iu/CWL/FIXmJxSo0vgNRXGn07
6XxXd1gYAQiIPlmxtRAr/SXY2khZnmn/wfDwmxU1MVPMENewXaHsjwaykX/cpbkL1iZriwUk1Qer
3BV8JTFKn0ac6brPM1nMc/gHYUfX59YZTZQ/rQ9gZMf7qwYMV8qLawQL8sEFWn4ZRNH5nxUNS411
YO9rNN9e8dn5UaNyu/YY9ceq1NeBhxh3dfpest1yz0fnqiwsMBeMCyjqmqabkfXUv3t72kGrKTtd
wSCRESe3eRas9rWEqiqdJKug5t3Px4FJHeLE39SXlAq+O0Nm3EvQ0fUOeFb+A+G2JRMYi27pF/+z
IR2FyxxHUup3Az/368ZcT4NmAVyk2IeyuNXThVuTP1qKfwAMgxCA6/FHQwG1Us2ma+syF5qIXX0f
zOFkaXAJi5vIpH3+95g3aLi/Vm9PHEgvKWxldhcUr3GW3QzwxrXlHEKrl/k9L4Zslu+lBVPcN0Cx
iruOxZUifOHmoNgjBLSdui2Qyy6vYYMUHhPBXowdp8i0dmn3peovLR83pgVc1r4YXQGxbcwh4F9o
JXFYFQVVn9rDcJpwvvR4DbFeaQKnYpYqPA9S46iUcCQqFr2BrM3tV20JUdK6LyYwUfPp2FiKY8Sl
nz0Ddc3i4DCqUneeuHUAoJ2freSggejwuRsodm2Zm4eCPc0M4Z1oQLUWsRFvCf0Y8hUfhlp+nYCj
niOv5ecjlQtXveuGU5WdW5WtZmOMRUKYsI987jj+QLlWBLfTRGdbToMTJQ9Y7r+f85Yntqv2Vr6q
EXjZeZme4OJVh2GDISDjH5lU0pThnfKQyLXJZ6wVT9UQuHOlGEcTaWEFZrZtw7NhDmO8Rrcw82Rk
EHL/N/WH/d5E+hYIYX+s8N5dxHXNzD6Uz5ab9jDfsLaLuoEvszYXQDudBo/+jU9SaNVUEbClExrT
n/J/PKXDExs6/TbscYdsG7HRxiOAS57x6nmJmA+/moySTlbdKkqnQeTw9Mp+ApTU+l2a6aWU+LfP
bZrjqWSRkBNPOqHA4uixbV8WX7n7dqH4FwDn3zGGORgfy1+6kGA//7EhSVC6HG1e8g0+z53ygAfj
UNMk/A4DCiCXV+QTY0RfMedNEcg5LxBGj16e+IqWwpMrXksB/lF9rzXb6X53VrtKlMkJP8q94P8Y
pTiQ3ovw87rVCtq4CWtrZUx9OzquhU/sZF5ih2x0lVrvyAI/3ixe4TNqGo8bKHWB324qOy32KjFX
qXS6cdilLNDkdSo2HsWj0sMuPY3mJ4s56sC3ic63tgL6bRpQY06So9KnO0ZcQcSDAs/0wqKvnhnC
tbGzqmqtb/dfHEXA56rq/Y8KIrwUXreD5vSBlI11rvh4X79b4vzW7obfoEhPqCXL6qeJ5q6ad2AS
6P0kKg2BR4af/p5c+2Wbk9eWS44ekllTrKlHXA3XuKLhrABB6UoFQnYXJUr/XKu+y9XWc62X8vCF
ykcpyNMOi8zl91g2555YcBAf9VrpIAOh/tdPf+AhxHiYfQo9W5kiWCnEegOjk2XWUp1wW0UEE40j
4y7V+E3CotDitKW7vDNCTpCa5fkh9ZretG+24fhG44Zd5yfsz1RtJCgOq5wZdla0BT4su0RxWUJ2
YoVoDQ7PpoNtoFbB8RT1b+7yA2yUvxXphQHH2LPjPkELezCj4/k8bxt6pxjyM8Vz21h7UwoeZRWu
0+CzZ9crLhN4xjXdQC87jibpvLN88Xaf9VukJPxwlbos5KuD0qrNWD97GRqlSAOKt/OZFvUzNKnq
dxQVAnMH0MM6xqR8awidAD5MgbwpYv8Y6jAQJKRecW3DWzMnBL9ANUcX5LYN6EmZsd3Uecbag62E
D+9RFf1jEN1Q2hTPxRPJe3C2SzEKHfNniifdtcuGnmtGbLHf5dWdRvBdhLMtY79WklhYYRtHVAr+
X/qXKf+XCxu5T7UIJEZG+iV9v2RSixDW+Ubmn4kaL1vVt4ksgGFa2Z0ki65ZM6dYr3MOFsZqI6E5
AOM55Aqn3E5OqK8TNay/VQkC7nAO7eEFH6Z6MOtF2QGJg1YdT1ky7XRwHzmoWdqZ0KxYaA6IHNqD
9lYcQ+tq6hm6oCrVpiNhwmPUyC5sW1RrFNwTZP1rT7GdAlxS+T9zMdXsrBmrwUeeI2t0+l0rhzrn
0lOm8Y3OpD4gbkDgiLh+pNGwfNVuODn1nImdGorCqrzVhNXUu/dRGpz3raE9pfmMoFoLbcYQtkao
LQXMB9RHkguKYKEIOachReP6+Yunprt731JD5FYfWS0z7RegZy/nxphxv4tzAnSCGdcZyLn8xS1W
+8ShMjuOs33U9r0qnr12PcSlw7S+H2ul9dEKlmer0S+nfP6MEkiAQy2sNCzbX5RkV6nhWHgktuMZ
JrYMuXCxUv9w7IN5eSCSInV0N2YFE5VCXSlAPsqXAMjgCOcr2lMEn2zjIqHfqNSeZp2qPXscGZ/e
Ur1+MaHJhJQmXIavboYhZNXDR+7PArqz4lfIvSr4eBy1rd44XtVbjE6u5fbcma/Fa5k74AME1OJ2
AWtUQEKCs+t6/pcM5R5NrNeqfokLfEfyDy7p0w0k7J5QMpUznhlqWgV+sy3kVhkVMuzeWxHDPY7j
DcE2QyAO/txCYtSqEKkOqjZG2Uvm/ASvH7BgkvBZcLRlyJ9xfafYcNWDHSMT7+FYlZp6+7TKaGvD
oRjokPKYH5zI5AMJgrrv3nhHrbGaYumtU0W6KGUlpqKVXcyhxTNWqQLfpjXoGnoK75YLTUryceTq
nwmnf2azADVpD4FA+N1V4ISqzoMXBPMH5J16T2uTX0FG0iH/sys9af6L/cPIYAMQvDyBr3DEm62n
iVCbah/vp+nISUcwaxSHjb6bP+K5RmQ+Hl90324WzStSJjNNSzBFUO3NP3/oEIhds52U8+q5eZSd
n5VWwjTOvmd5hdkIC/dYZuc6JYuwUsC2jeMM6HO0RFUsAJrn1jagykecILFEkv0641I/KH3Ldv2z
qwZvQosgd5YP/Wyp1iVfH7TFZ+8g2aLOlWXxXoMNZsEKxKO2tHKvmTshUkb4anOxKTv4oyLCAaa0
F8fTaije4SdgNo5cgZ5u++uTeneSxGAZAyyESl0nKhQ0fFA7sZd4oXWu/xLznLO9+iCHr2xiP2i8
lIUc0Th1xBTmPcvKOqUCaczoRHwZblFIzE4Kn6MyZsle46NZLjct8dPr9iIhr13wB5Oi63xtlgdZ
5mFn6U44pP+j26pX8K03PhXUVF3JdyxYwTRqdUMQ3UgpwvrddG13+8vkIgbXA5zj1nEQicIDUQiC
lTAWRlUHzo16goFdhtn8FpPqu7WGAoKQTStXpJ3I2gtvbfNtAokhlPeU+910S92Y/BUbwEQIXpOO
XcOugMivdBxX7/pHmFatcaNymZaJaRik4a8EmvJUvTK03LF2CuRPi/QZviouN+6v7X/S8oGan1wJ
R7vCGnj+2jwxQa9X6TNg6JJ9NFQUkSsLoUv07XvYY5W2mYyly8UcfLKDStm3tpAN/0ps/6LpUqE3
tq8CskR5EF4tbP8tU0lGAjk0tB3fK/sup061twVLcbzZLyCirbTlrF95sTdMFwY0+EEmv+B5De49
KuiUIDu3B1WR/bB8nTHEsFGtJ99L3ziRA3E/XYCpOUDiiAiEllnTmDqbfDwxXZ5aXFIwJl4dwJfR
fBs7jB1x6Y3wbgqaKA9GTMDwnleRARpu3nqRxSbgHZse5Sx9QrP0Oq8LT5+2r9WceEcDmu18XYzB
ISCVJMcSpu63YJXiUSTswS01eH+0kwqrwlIWBEw8sXZHipUDtBIDD/YWcDM3oI9jAeh4woyBLFNu
1RZ1FJ+X0uOMre+zH8Ug3TRkWpUFB7odfTIxeQBUce7Y4NW5Ey6N81MQsQFvwVHo4QggeVltA7Bp
XfnPRIc3n6HuCKI6PtV4c7UncOZMQadP+C14GZDo+ZeR64hRrxwpCRs3+g8h5NNKdh3u3LGEDY72
gIJuDX4orO1OKe4Or8ZNbXE5M/PojVX/ATa5X0YtdI32TMPD5gsPeK7TuOj0TZYqIf/mN4yw0xwo
vaOt+AjpHaqlHOSdGBld2rkYRCZgq5unF9/sDOQcvYAYrdyb8tlzVhalg1kNgLe5zxImKXz6dPhh
UQUct/so7/bXwX07uWD8TZ+o+/dCdCU9LG8WwjymH5FBmvYjtiPP7VZdy42lgPbyyoq7NjTBDiyx
HEDX2zwEpLap0y8ihvc7/7snZJ7krOpWLtc95PuS+Bw7vuPPzmbl6c8FE2zU3oPKq+G70wTq+aoh
HdYAHNFBMiCu7TC7VlLjKZ9jl01Q/2unUpQYjqxJILdUMCYS9tF+tdTppGGCYlIUvFzW/mbbfl8+
q4r88DLCy3BgvcR2+CPawQpOGdg8xvrEGURCKBYsG3VNCAdJBYTPifMpYKjTYZRxGY8GzapMhYOO
J0Pf2p+jfdPs/oQNs78FR1jR41HVEP0sD6EiFWWK4QnSDHci2CMNVRHKARge0HxlCtrhAQJRvNH4
AO/0QacmmwUFB2EO40qncij0Yg7xW651aWFr8+bnpMjUAq92CshOoO6fetqAXkrRHSZpmTRf0nBT
Jaa85PVBCsxcDO2rXyriFFDyju3BDb74+Qbn/mZyfU8rAt/mAYUCiw1U01I6AIKEGAwK0IcjV3OU
uxY29n4fBjd7kogO1V1q6JjAbbEJ2wOO011aLciU7uCEnbDQ13k72ImlwzgtpIgFm8bFQ59wQjx+
j8JI+YKWKMx4mgHmHcFZbTU7+W9vj1jFtbU+z4KiB+hi+4pXa5g95Gt2mcF6jFqarRNGTosaJIsY
SjNafh9yGJGJqZocmYygwXlkUrgjXHzSJ3wD2Ee/X6X2dPsSts5xLRcpDWVGgzkHiTXymCPq/aFG
QmiERvi2QtomkDHZt5SH37aPdGTZKauOCN5xmW30EypWQh4Sua3wzVfUOExgsQiWLIlKeJUpTA9w
6uwoVPaK52Z4b/aAnjP3c8ccsXjHHHBVuZMJs0/R+HgLUVUKXcAMSsGBgjTc0mcgYTN+1qdMwHMr
K6sXgbpaBkLmSdYJR6mvBiZLB8zwT88LjNQxGYuYys8kz/+RyJjZKq01h7S59GBGcbMRYrprm5SV
/2efGCgJwCmS6TJj1o7wlO9OXYBM/OTSnmTrPSxl1qlbuh7DsnVd5hiD0K7TpTvEJcaDed2P4vMj
CR3HTAIxMD2hh3hKMoBlKGY3z/Pi8yFa0qVZXAMDJXX23rx3r1FkI5Sa1HPAYCF+Fmta7am8eISE
K9An9wh/oHBS96oIbODRtYo5szj87J7iB1Rqme1iGK06s+r/ZXRDB8KaCgqIMJzWh3CfTGxRw65r
tXH+ZytvsFHBI7cjwM8B+QFmzevVnADXWMxtRCl+uRP1R1HJI1noBGwHYnLndQFi+0QVTw+xv8ig
aCMLa/5qVa7MhbkoI3/MwGZsCzBNUJEwj6CiCy4m9N+bqfruMVg4kxls02iUkOqm/iwhmT8s0UC/
EGodoi9gNbw20P2+av8h+wTYD4OU6SIYRERNOsNY1LN55xnDPUoUZq1B/nkTuwe1Send6ocXojEa
XLbDw6saNtDmHyEdtD0LVzmGzf+wmACyanRnjwFItGno/mhg2sZYJzyyiG9lNUhG1EdsW8aRigUj
bPcmnGsuYMZvlmkYfYhLPEjlEz6NQ8OmbJS0XSdkEsumdoZaXT+DqwrPYETh3d6w/MxA82F2CyJJ
sWmMTgByH26x3KtU041qqlvUutOlRaFinacQz8WBN3Wlhp5k7Kkm03Z/Q5Ls7PHVhn1NnIGicoTZ
+60/TlnM8vafV6GQdJkyvfI5J/LvVnFrsovEYf9MN9zdIaaOqgplNCzg9zVDoMVfYLtLzQJujCtZ
5bGs0X9CmAt0BnrT2EA7gM8faLkvr8dcqSl1uDBbj6Cm1KByeWqOwuXxys0rTI7djpUPzFQpAjUO
nWv+6ItCvHuaT1SKeL4SNMQCG/a8B6MlLtZPnaVv4E2bQUEQqYyVSnaG7/FWas9YuSeLgCY3AfUh
pXu+Oo2TphWTAGpT5bSt+QoAEXv8usKZIRIltlElRDUuQ18kcTEZdAaJ1pvDupojyB4BQaApdSAC
tR3W2hxVl/I4xh6J9OUsMp58ei6ayq+6FB0y/PvlLXZbkLrl17AIjinxOVlF5/qEODdD5Wvo/Lh1
AGDZKuu78SnqdnmyB2zGTR2MH3EaYVLCnZTHTUu0MtAOSuHo37B66e7BBH0gLfF/4DgaD4F/iaM3
8+c3QYo7/P5VWDDxfayhT+XF7pOYGUwGxmUuCA6nOqVO8QUSuCvX7rwWA0FBUh9EWoGfDSXah3v7
syXbLqtqwAN7Xl7kssDg35nOGKJJvZ5H42Z62ptLrJcYvwuPwI56syYrQ0WvV6cHvLEPZsBqhz1e
dmEaGzQbbauhgtg8syJvuVYccw+EYjH0A9WVc9BiEsRC0VIhSI5olFR5kik9iOqXHymhEwrHCeic
NJE2MRJFz4TzH+f7lxE191RghtWZxK2z5+r2QnYfX75s8iKZ/jDhITWJp4OpzW/qFBdz1cILl+7L
U4la7pD59MIgiMqkTPk28Kh/bnfIGZWj4iVPHdrr7u7Sjc31ixYCNZDvqzF2nDYCoxYhTwWEIRcI
8NoFpjod71BK7qw2wm0a8HDKCNVcUbDu71ktujJA65DxE1UJPIamk1IWORYVdpXNAdte+wmz27n+
yP5BMF809sMi7K5AR2k95xuxu7ElDE4Z5MHnQp4blFe31/+IJtiFspiQD0DXVbGuGBgwXb45yYBx
R9VsIaN/t/mZ4B8DeQxpOrN5hA17Ej0YXeYJrfYpT1u1iiQtcLudYVhQgYhKGQ/7YlaZoZQw4z8J
22BjGxDEx6/u9jHbP6UuXlfLOAOfHofMx9szLE9Z/Bu2w2lMhQgOdB1rgn9MbJ/YJBjyV7axgHB7
BUE6whNzEhJKrW4z/6aHwVmxQBJUwPHiDjMBMGeBQS+J116m3QhDwKq9aT94vNsduJvOQMtLAIog
damlIZlHAJAEf5M0c4F1X2q9aSRDLGmGTTyP6PADhjXyey4/3ZBRTsToBgd/hPuPEcknmfCyzQZx
z5JDsJ2BCrZWtIymnV5+PBsBctyhfkx1l2eLSrDc5mdNw7pi6Rv0YTbl+chuIBKd5xxRuXbCbTSZ
Jnv6E5+rVI/aFcIDz276q4sy/OdJQj9w7iUAePVvIb65fxjiElIClqOT+/9So5hVGBE+ZVBDGV0l
8qbLnavQA5awGe8JH7DFgukxeicXPMISazud0oIqmlh8Z2rrnqxskeaJ7/szf0MPBj8C2GIItv/k
Yg/XMaHY2K/Zr29a/AQ6+KOteMZRIpzp+G5CRzRXk0PwCctYKctlnVarYwJkdcgi7a7TPXhD33Z2
OEMKxc6GDwwEusPhsiv3bAffM8+IKa1mtU5BKGuB+BmXJBlIs9nZUNtcU5nu2Fa9SBDX0Tqsr2wK
F6odgkP31g5488Byjsi4mwzDjUJIjOgLZAwxmSl5CWtxXX5gjWG0mA6PsU8Xl5dscLNEi3lgCaEh
ZnNdQLt3wMb1WUgWBanEmgQwYTC5i93GI0tdrwI+uUA5/sJL6n0kaHjyRdsaUSUYd/7Qsh5Qu+t5
ACyDLBg49VYuwL4FRfxkKwwwCa8oq1UibthIVPaAErqFNhj0trBwAKo468YYfohZlDdI8QwNCE2o
Ehxr2rJR+YtWWsq3rvBv3Ou81jDz2wUyHVKWQh/Z6qeRtf1Zx5S2U2XGvAO7WClt8hgxOEBGljdf
Vucix0Zm6bDe+5qbQwb5IlrRCBWiotpnODQFHQLzSE4mnASecDl9GQ3YNICrUkIxCELzvDB+GMfC
PFgf4WZY46I1Hvba+Gvq7aGqMatzNHYdNMpx0a46F20P7JITxgwYjF5+sNLM1DwEKp4cD1gdfIqc
Uoqr+CtQrfmrreXpD7ByvXf1Yc0ivcboEBO9lsCaL7j7lkx9qb09mHC9mq1pt/uayGK4mLbX3AZd
Njhwf56QtyLWfY1wFPs0PozzVWTcxXAqdUgqMScowfON/N15xKlhznmzkafueEN7ii/U+ezVHJJZ
ZFnnCWbKLZe0Iv08WjE0T+vrlR8UMyCpDlZh657utQTsdukECo6wtX31c3oIG9/vKHoJlFZxm+ns
ZGbr4yeoHlpESSrnt/d3Qdr9PkTP0ZWQNTR+gwGU2lYVz4e6/s7g8gb/i9FXJauf/hJNjT6CMEPg
iI8GPW7GRNHGjr7Xy6834e9vusM/J9ocEVmVtrNyo60hzYNwczMNTb5KncmIOma6Mn8MFMzK/Bdc
h0VnYNmP/eO8lMGMnS9SUAP/IBVZl7AFnKnk21nxeVWyEmgT5TvkAnT0JhVqRZM8mVpr8atXXx5x
YgPBNMk/G6MLFQc9Tm+Ts/PUtEw7wNsIoDu+/0Uo+He2t2+UupfPxL9M143MB9nrDVi8KUXh9dDm
2QE0nC+W2/817T7riZnTuddQozCG8rabfr4tuQtoUqez3JKDhgol660MELjC+LxPBSk2dfVd226K
y//0yLmrRZWCnYJNW/RSXzLrt3azvHH38KasYr/Yot03XN3eCbHsepcEx38NLwodUTLJ/kp68V7u
9qUROn/Z5BNKdN+ihCSsQOPj6QyzJqnQCNfwb3QKwnm1/hNvNOSTFkm5r6MJQ4lnHaTftUfm508n
vu9LueXrKvyHNGtI2GdxWdTCrTbzzUj17Wld2DIAwEgGVqGLEtCpXn2DR8mKHatAia2fSsCplMkK
zch0BtkP9NzFWeMJM9LKovYeRH1Yrt4MEUo8zKrMDegbjApkw020tSWLeU172mWm3zGApsaiBiU0
CnblqdBKvmtq5qqHdRJOsZCn8DRwjgEROPIRYWzGjvEOsmG8COhpI3Niq1lSufOQphYCIuL9DV8o
NAJX+z4IJJToJMLSbQ9Oq6C9cz/j5VfxVBVqXaRPav99L4PqF8GQS5ofB7mCaoGkWmDvHPLm0Biw
6wYvbCGaOs9qHMC1ywgb5PPE7QVykbsMLP7htLBEOWqvm+WUZMBNSGpPXnzG09KZDmHayDN8fWFH
4y+EM8EDcEt6kXKICpkp0lDs8CpiO9dMla7HiMbXMNzH7jpXM0YgcoKTW6yPTe5/gLP7qhV+xO1S
YFvqTJpogZg/9a2Xw8ck79Z4D2lguvp4MuVlTW9CXicDTv3bF1PR2BlLp5iZyg7AVYluEV0ejzR/
3hmcGT8HipFttMRjS6y3VXZIGWvSe7edtXp3G7eCTwy+dEQONXOlDlK84/zTBa6tB+invQb9cIZN
1ifDFeAFCYkQU8/ZwcaRWfmtoPjvuLeGjd5rzbmV5qd/0VpcIBXxSQy6YhH0tQkCeJo6I5nd6qhQ
YCixTr61mBo5ONJ8TPeYmNN5oXWqONqG15GgV1TLNFoDF7RQabbPUMh/VS2bawWtgtp7c5jjSZfF
ZhOsXPEpDbaR7J5R6Fe0lDaWirggH3zAOBb7C1Hvr3c8gHUUi6h9VMpAmV4qfKt5AbVHRhYsqxwK
pkNImrgjQKgXtvP8T2ceUHXlsd/CouOMfee4iUMn8yM81dkgDl4gh6LaHpvu3eVK4nfqIByKQlR8
9MuKdPmbRNQwGr/xLzgPibU5hDQKFcOtGI6a5I8kXkCjpa5XOYiChDLedy3MOXqICu3HoletK2V9
TW5uhelDrUuhxP0C/bU3ej2pfKzKTUBb5wRRzlMpQvYy+HiL31VVwYYBm+o4J0uQs3ADX97+vJlP
OApVqOf/xCQkvfPS0cXG0SmsC60FddnulOFZnJqMok8MBUNSFiA3OHkAgKIPyLtPDoshUtWNUV0h
W7oOZwx7n1EL3nPurrNhHYV0db1lWxU6l9yBnjC/O5I3MfDpLDPUkx0ORVRYVL0oCdrHzl2Ug9Rx
Wy3V91E+289KtSjDytARcJNw+/9P7GMKw8mVjO5qGBei6YR128C0v0uhej80wY2SRcnz7twjC86v
w5D4wSDsZkCvZDRMsQ4sOIDI7BTICjD0wSBU8NWxURdorU9uspGijnqYJ7miKfuAWBVSctKYfZbr
/1PmbbJtCnPSwrlUHW+NJmE43be5Ku8gOR75GInCyuTVIXYyMZu2gXtOGQ6GKhvAuwyVVYVswbi7
9AyKuIhCnrzvSR7qhUgn8aRL3BR/eHD6RnrVAD8E071McU5bv4o0wZp3XxZ26r5ucAwVc3265uGp
ki0YyFii3fB59nm3MRTrGT7nDse+v1bqQgOzlnwuzujfy/c07rNsUo2gl7sgARra6F2Cr2p1NsWG
+KeMa+zxYpzl5eIjglXOYszHw7ikvwolmsy/x7xjHu03TzoAhe/TU3zHbNMYuUbSl6qSvfTFJpH6
aWETV2QvAUqDz9VjqeWOpwpp5sgkse2t64Pj/reS2TKTgql1wIUpqEr4BFjnGN98E6lB5K3mn7j4
U8ejYA2NdoM9SuIjwPqHTgvwAEAFMPwt9Hanz3NZCCPVrfPGoehQyt/Mkv2vvb4afpvaOIvKeLWo
SSfFjVjB7xKRrqD9s9ZjHuVeBgJGc6QSkqJQJP8rHsKCzKCQWnsVZrvwcjVl4D2z626qUUaFTa9d
DMSWoIlqAPoCxX2TCz/Ler0A8n36vqilDd8WhVZKRGokltTUaFfotDb+VsGCX75+fXA16LjOHmVI
v6q3FspUSkoY/S+JovsPj7EDe9/f1aMS/ii2g7M5pXkmQ2M/7k8Ur7gdtAj6AYPljAUFV8LM9OyV
V/JBRr0CVMcwvGkB9GQDXb4zPFY+n+B2c8uZjXUU6NDKuNfOechNtiGSB3xjb5PoI7UlXHk7rdFl
RUdytIyoihlpXpjaMrh639RmLhXqe5joeYSI6J7ORSImrXn/USA6q0BMrKkMnRlgjYhLP34oYDGv
DT7QkWIM7504Pfh9TK7WNJ2ZGTouXJbpGxF+8WgD7mwzYwOqgTvGAqNfenlX6xwjHqItcIsti2dK
nxFysU3bokLyAXKqdiiSzgUuYUeIwBtEnx10W8XDMIgWAVWje+mI3qPnhilc+RVodhL0YUUsGmeO
cGSH9g6VnZsmBtiqfwvMULoqfzlLveKKHy1z1cCP7yT9V5LNhoq2grFQSwMC+yLRE+KlF1O2lA2m
QxGLTolMp65rIdA7oeeK3g5y+hvr9hauI8wwvUnpHnrKFSI/KE22rFdv2pJ6rHwDKD09Dt+cZqmM
c/CJXG9MTf6dxVXxgPsyZFi1BaITv0hqmtlg7A6oKtU6blMBvjK46A8d7H5cPN6u4M8eWsKYQtpb
tyteRRuHBSYGsQBzI1Cy0VkoV9io7HU9IZ8+emjw9cby1TJVKGgd2QdLR/UnQSJeNtRAyRCg2w/2
7naVn3LQV7PTK1AP7qY1hLUsd8IeahejPqy851GC4zo8OnRTHzhG8PrU3w55xjZRuMhuXqsIMuSG
AhRWzOXq+04X2fxCO+6OqUrIFUGSvljpSJ0O0+Y8w7rJE/+5octtQKuAvnTJO5AwhUHNNiGvhVfk
wvVEfLvPl/0JzT4uk244sn9egQsUIif5yKjFHEaYz9DhSng8NuSwgnRt/vGUcH+ztFua1TXQV/8T
fpobpvZYKdzn5r5tBDPVy2DHM502M1eN1iV/Nh2loCWTkq4f9apJg5L2WWyTSbw3PJxYVM+YVeEK
ST7ttF9e1z2c4Yw0nIf4rNICEms1J7CA6747tJEF7YeX1KkQ0leEdt9qe0CdG1DeonMIMqWm2xJ1
rLF9qkHa0A1XaAhLjZ2keDt1NLbYA/8QDcZ7INvyeT53oLiqkwXmtJHLkmHYu13xnA1/+5JgZg9z
LmYpe+i0pzotz7RJB18sUtBkgJ+YXTkdS1Cp/rUwnR3CYKFV3sk+Ykla9Uyvc6iFzMlhQHh4Xs39
CVxbyBs3qoTQ9zxTb50nA0mnmmaJk+ACON/vm5yqbcjN0M80ftp2qDQ+4OmVYrZLdX5p4hQD+ZeX
77oPYMReCPvzmadznf5q5hUZk2+ylCny14+dMAKunQUtP7XHXQCMxAMP2BGl3p/SlQpl9eHNygXe
rVArn+KCmgnbBV0RMFZaqZj4wsFGnbv2dXcyVNIVta57GLGoV+8LRFC8HaYG5Wyl4DMdUEbT2XhS
U4r0UXjC2xls13A8EeTKAT5wOywLXdQwtMUw+amHbp7zkC1pxtF+pBUmBvrIEL2KVPj+HmYWLX99
fH+eMC/JNuv/+vnHnTkEHc4+p33AoN8rPVYE7wdf4fhdOGVdMzFLCmIKacM52svwcuxbx5+PPc2r
+UuTLgwJnOvgsRnKrjWu2i+iF7wUa0cBfio7T9kYmAsJwRjvW6dsFSNJet7pnPM4iIdsFcDQ6hlR
vKZHE7nLSw0J7dy9VaUSS97ICFN6AZkQkmSMvtzFHIcLpNN8asvujjwYomp+hAr3ZvwXvtG/iRN5
2voM2epvXthNqAGEVIU6Xkq/HEFdmQGyY7D/+DwW2W8qaa9UNk8HUoyjkJZ/Ps3AYbSzRQ9SwGX9
0iEBCxd0RknTW5PwaevKurRbwadc9LVv/M3pWJfpTPdwAJBsKcHPfRi/g8uibaEBaVmpAdsUx4IN
FN5Rp4s3t70lhw22ww8vNveTlRRshJC43tiZ7MUJZVKnuuyR+8PUG7bNX68UwhhG+DjTUqqU5+Ef
x9YuRz99BPZxw0OOpuPnW5qtvpE71pKz5OxrpHm/+Irjf1yyxsmiLnAUYbKXqIHHex+oMK1pN1Cx
7zc63kJCl9Vu20Ob+aX5dBNl2mV5oeZFaewRHKnzu2Du6RME7ZgszrodDG5jBpXW78kn+7vsR4WJ
ZyuSkCntKl1ZrIBJnekxPuvy03Yxnqs0jobhO3UOdLZzEPilUwXv/DBS8OYaJxGi7EbVQBEKbZNF
VfXzSC1QzAwbMxPV5GzCQanWJNo4VNZg1VNkdZ00GjZBr+r3bYOC1z+di/kvCVYDKCnBp4fx2/af
8zH8YOmCpwlG4pPYYf0qOmQ86mawmvrdFyFEcacaaqVIcMZbFYyfuFyiclaoJ4qh87jYFPwv7uxF
oz3EtfArbrgWK2hKlTQ6BE7Prjp6w+hKa5rzr33Bi9dnir0SJiaN0Adkd9V50MfC1VkygmMBMnlO
isPSXaQElWWwMWshqtKLfEuUwHVyhCI8IDO9FzlusyApTicdFYMKjBJBHkB3AQ6FRPJSbiwWHpBR
56FHICiv1QccjHL6EGQm8TNXJ2h9CYqJHm4ZYeuF5H1HsHTFjM649gzoUOQR/gDFhg+QmwmKLeKv
Dhk00zOTSoH+dvXzLMuy+vuMk72tqEXBWw4jOZtvASOXKLtrW6T9BYUFU83qCNETSXxeolAJBLDW
xQCHEcUQS1MCClTbkYu4+mHgwT18zaIINuGr43wgVshJDzK0KVNV6UyW/sRrfkyGV3He4H2kN51D
y3VB7xngMRg4SGmxN+cuChTaQsroT93awft+UpGta8W+F5/nf5n7qyqgNxoeYPWIbMMamSr4+jFL
kTXWZf+S68jz48nh7n1jceQYOOpVgSF+ZgpVp2f+mo0KHYhQmX2VZXH/N89iOda9ulYO8y6C5ni7
ZkE3apCaHveUofiZpfyq1No6+XMGe7NjqplE9OxaovVfJv4SH89sI7ZfWSaOmQ24bsElJDO2KVVs
X+ha9pxONHACrsnnG/nL9F34OIa0S9ObKqUHM8kF+dA8c7sJVfEDpzfFrFuVSq9jmXjFWOLwiuEL
kx/19wL9XAwJxp+L89A/gGofXpz9S2H1+L5auAxH4rT9DzF3PyOyma6hN+zVJuiGwWbocrYvxtwE
Fs0g0lWzifsFx3SZagC77idgISO1jqMkRTj4ZCPnPT8NVg5MhBTtGv/t4gOZi9iGnJGTCPoNsLRt
V0ndZVLXC+Ia3J0h0u3wS0+mQM4NmHryPLdpmog49dVBY3EBtEItXMh/wRjjdbtu5ZWClrXvLL84
+fHxJjx1OH1H3XDGlV9rhRzK2F7Gyk15ecoiuOAqXX8/Xn7FsJjsGa5GtpUn9lDOSw+3Y6lYfzc8
0h6w1iZxsWRbMamjV1T/DMLD+OnW0B/K0S1/r9Op26Xb3TvYMvbSf4e99Y6z93mkT7ARpAqeAFgA
IZOk6pD1hwRvg4n1uCY1n1AxZDVvKTJ3F42XNYL6IzZurCpcJO9azHeBKsGNr2Z6etqLfYL9u5a8
B2aVNg58sh+ia40B0ZBdWe/A1Vfa+ekZbLXqYXa4XANC3qD/PZtHFDWWWp0XXH+xzVQs8nNw52NA
mLWZNToOth/hwLY7DeCgFJUtQ7qfrtyrSHpjy+QCGfTbMERjxePMrlgWovrT7fNBZgOxhiMIeNme
iBWMOE+lysoDx90VzyLd2h9TSkSy/gTdSg9osPfiE3t8Y76kQL5uKZA2sY6Fbi2s7J+Cos+730ro
upZyBEFvdn/hlR7s9L4Yl56oPtwsleoWAwJG7P1X66myprProSEtEj67Jm+HAx1Py7wcBwlM24FZ
SgWwGnRMNMsusgcK0Ap0nSFLu7Vaw/bwbyLQQKLYmMh6TMpSA4uqAyBlSf3YxoNFiVYPFYCO+WeR
fNQ8r8cNAyK7cFweiNmitJknxc6o0XMPhxuX/Y7KKVoKAvk5ZKbFtmzu7+f0mgFv9cSdRQyTZSJO
fkqoLuG50NshdPIooQbCslixWEbrYO2xzXAkGNT/puSrQoAkHqqu8LEC2TuI4+Gsalha/22DyCwi
evcEzu6a2PnhyJTX7/kojoPZn433QLt7NDaE5NB6sDrUlCtQ7FKxF/uM8nBbmEsa/4LiLagP1TBK
a1Q/gjOTIRvHKLSYlW5poQdvlfq4mq4ex1akPSUGcoVFurAVnH9EhqyOdHW0tpTfrZMhkUDOnrJ8
nhWRW7GRLVsV+PLcfPT3VJL7BLMCKNAnUnTOUdxgiIe4sFrFwGcomKJjJOz6vpp0L0ZVi2DOZv+n
T+4gLKbQKGHYWTwwFygpm0x5W5qAjFnWaQjhf52SpjD/OsdjDvWxjtC8MYlsQVt7W77EBKttnkMH
v4xE1o2P5fGh1oOgxYgaAdQUlyTCkX/QeBKqJIsVyBnNKKMtqJGdlbYt+nXTjpqszURa/VPaFNu5
uDg4UsxsZfHMuvLADMwbsEka3jdZvFGbbfyyw4qcYvwLiVRD2MHEaGTREjO3AZqU2u/3Jy11ALhP
vu9gspZenE2CQcXAmc5dFgUUup6RKHMzms/DHhjCG7a4yOP5/11HLFwiKmp6gQa+D3d7niAk3zeL
oZO/nkIS/7AqXgXk8QlpBmlWsCyUhcdoK+ywyVfaQd5wfMhDU1vCa9BD7GhsNo8I1VZUFjPhiiEe
7GzUKqS9+FSXgZEwC7wbHLdvYRADyOHRnjhF8/Vm03aDBlAYXg+ObUMoxQ559rjKNe0I+B0uNTQo
rm5QcozLn5R9MFQlg7g7klTyoAvuwmZvGFZ5lrYlWZ/GDif9V1joWPdcUrRDtQqhfol3vOy+6OSN
QZCvaCjlCg4f15QoQHqbzjc3dj0UcC4ktTJ2FfksM9YLw3RVBcZLW+/E3JGR35HNMA0pAYHf9fSP
8m0gAVHQbdHBWvBiE1HBE8Rs4lqwYGoD72hLVJNEl850fXo5OU5eyepPjDAd3tGipPCsZKecX7aj
TcrlsQKHU5kQBhmCJhkFTKahGYPL/RBw0HBeatld88IuUEurZvNIG80BeOmO0C6PCE6Lkb2GI9cZ
AEsXBY3lWaqrycU3kqZGQiL1PiY7GJPGe/1Rl0Hnm+Dzu6ICzQG+5lUWXZBP0PxbEGs+eV8aCgiy
nKIWi0pIkrxSMI5PC7yAHirEil1ofQpmpDS18Ln1xolm1XtalTqsaOKiykdQotRrTf2fOJACysNL
Pi/Fj7GZ2D4x8ChvfvHE3qqbF/IMlRIcrW6wyuWpZxFD6PKqAZ7+UVeZBjSAfEdiyvN0gr5w8u95
TOFZqeLPvmg6qLq5vusj4PODNJo2cILHraBHq0i2VA0aJK/RTcNUBQpQP+x3xwHxdYpRTeBK9Q68
YBQHXwReS6H0PKZD0x80wsh8PSuWXJQRT1wKTqh6fwNhBwlgc+qHiwzQC0hOnaDwtXbdL4Tv122Q
J8PGhYnPeKFaj53wmZbO8FNb2TEZ9ZhPx7ixyCEh54tWc3qIwZ9oQkSBKXOOxi2xOF4Xyp9INWr3
8lET2HpmZBp7JrX/GrAJuUFhHM50GGhuDismfeTcAQU0tOVq6EElGwfWl7DmWR7fL03skoV97cB4
PH0cBbzVwIM4jRLJe3BmwnJTwL4lTVFlHiWnU3/i5Kd2s1VAmE00fZDstmCStHMwpsWQyEdY4kFD
8xOcTLiIafJs0vHk7OJhJYY7FQIpJga7+Kdu3hZ6yiEgzpUUC9H/ysiGHdZx/WZT3zvFMvyHnARt
6lAUW7fAjyVMD4zNBwsG9pXp5KleqpREzTohfl7gteOW58Oz7N+gNgmCVzVWWyDNJ0cFXGuUtn6i
qFEMkAvrf2nOfYXXompMwN6etBdpj2ikA85WwHWVlB+6CerMUzJg4fbDl6qoAS95SiSxwD+RiS1b
s4NT52mrCeQkMSRl6lpk/zZxtqenIKSsWtjF7/XAAoAOKva0fgxhZ7qmUvZr2CLNJbooky0hHM5h
kleysgvilToQ4Sr+x75KUQpQHuLFt5kYYV5Utqn9PbZxM9k1Onn+1qF2L4x6z1+8YV4l426KYjxV
rlBE9DcICcT8ZHcrhJQcVJJQvbXo59e4YeGxhhvA3S0beDRpu4zlWkCRxlKCcRaRxlyyls8VnT2t
Qd7YnkDoksRhsIwPSaTB311q3B4RQas+rO7dUFZp1Ic2064OfIjHQXYJXt7RKGqUojDl+2mcd8dN
0ou0fSbaLW5tsSD4KxiqLRTpzHS7M+O7Rymm7OqaJlEhlRxY3egC+JGw3J9vcwLRzqarn/qqB/Ko
HgOtUu4OpVmK9E1ktxmGibz+gAzZpJ8o0a0exdoefKemzbZqQBPsnoV2jR26quc78BZiqzd4j4rE
Q2RE9ryz9lNsI+MeVbVy2DJvRmatvq1/8AFYXjrGZumMK/QbGuFYwV44T+DGI6rO9JOShGl3nlk9
1o59vajggVll/EMlebseOEnna2Nq/UUermyh0giiAkw8F4OgOS75jDjUJ8l+lhebRGH4kYUchUTF
0YuIWP8DZZGxJZmveG/vqggZ13VDeOBwlKnumBMJTH8pj3QFHTC1S0ey0sbdOUC9x4NCL6yfIcoc
OWkvUkJKOUmLghKUJY6CfSZl73b1h7jafYb5e+0EKBHUUXru1xNQ3idOw7HX3Rx0p/g3uvXciGAh
KbP0IPFsUUf/eROrqnggVnU5YQ8XziC6Vs+J/EGLUBWRlRdVx8+nIF0lLrrC1wZdxx+mZuST4SY2
8dgbYNGgUpUnjSOo4RxO9Vi4VfWhg7IgIT0xY+0NDRis+Lqawc0ALxynH3dDhyfofYDQ091SciER
dQd8CQ0PNpc/18LEls9A/cmbTLctFwGFHOuRbf8TuKIkKOlk2c5BoiI1YrJK9X1Ln5XRmmjicdu1
eSJaMrnJBKRBz7baaW/dDsBUIVC6Qnlp1h+N15iPPjgfnvYgivKMdZ8kerc311oYAoz4Kql1QKJ8
kQkqwZxHFztN+EJGXIdPoU6Rbm7+k9uAz1srQfJQKxacWsfRuLNJUfpwskbPJyZHPKS1u6yfDz+5
9+OV+wMEsQgSJAzs4/bwxqXmsZg+Lnrj8rmXGOfmM9Is9O9+D43maORVLr2EUzLtvRsVv+vzVWI/
k7g2HDiaMfyGg2J7rby0+paBbq/2UMkv4omOa8UAptG8ZLhtTx9r0jnhDd0Lr87qXBhPkOk/fPc4
sEMVKRw+P7iM78fO6DvGiBcD1ibZX/5mqjcuv0zF1/LDbEgm7wkqMQf1ikiTQpDMWOu2a8llMBZa
VfeJ0NLDnwedptpuA2Op7FqldsRmNvFbhmNfPSTAwd82zt2K1Ke1qXRlapQMH4cJXypxszs9EEit
4mL2PzeDFwvi/Bh6dph6dTSeHvWiULYutYZH1+a/EXGACd40AYh75QNjmVnHXOSfkc+qiXqjIH5c
B4XoDu5zkwGvRo2I5yziHo330QO04DH8bwfftJXDC898zlzLjHcf/IBoxtG/yxIvdY54WCFj1+N1
qsw4xQ8FmoOIg/OztTy7KZjuCAVMN50bELkab85+iYZpscmpNVPhJ4fdGBeALhpcViyWI6quSAPN
W/tQZ0Iu5OV+eMcpiV2OYUA4IwtsJJcJrn2lpEUoAQFa+jXcyXL3vxJlybGSmyc4ePK7j0ipT2qP
R8/L0bfzARh93QPmGRuJjxxlb29Y/BwNu8by6Y9yOljR85HTaMzQkXTGcvtg1afVHttHB2yggyLR
grhuKoSDI2a5XjuUAy9OPOMrKXmoYwQ4PjQ3fJ3rWt40DNCwgxCBc0dp/bJrMC49BmZHiDBUzZDp
dM1TdFlB/6vJZTJr8ypdHis2o2RE302ftOlNVzdvlHuezto485wG3WAyS+nGAbjt+xGmTx5156yK
aM5FBCMHcqZZBskHGDY/46wXEXpXXrPV354VecwRDZ9F00GC1magK2aDub0GAAfmK4vLVna5gXsW
4C3nhQ422I7J8fYiLM4OXdu25XOgG2yM3scPxEeCw04hS3u3S9O8wITxLmmlE2hitC9t7g0OR7g+
fkrlRE7BuS2iB0sVQY2O2hNtFxRoS8mcvfRNeau/fjKUXY5HcXoxbAEDsi9MiGntNyS7y84Ho3RQ
8EcIhOsebL0TZUmFbpuA0YoZVcqHTCDeliavgkGOszLK5oU/3r81FqYVyIMFm3QPzgdCTjajOQ5R
NBm2c1B8zWK5VXtIv63UKqmgvzpBwoPRbs4ptrt1Y8K6qblmiukKsXDqvsfGkd5Y717JgbHBeOBB
VPQTWNMC9ThbMKSybvfoPGN0k0Q3t7XUWDeG+puEH46teI5GskkLWrBIEJDLIKJ0YgrFYEQEy2XY
ViDCTbN8GeLjQi+ra5WRAASQwmtI3/vCW3Wn++4OP3olf6gg4aym4c8iu2LpgdqLFhRrKeb5jBgn
tctEKihE42D1nqQyFK1QDcc3l/fBmcpuSK4VdmvdQts1yYnLw0w26UEg+wZdtZ6MgxD6TjtE1cz2
8cB6UjNsojvrRPh5ByScW48tPMJjuM1sDSTo+HoN3V2eKWWrdVw6dryUCp0s5LeONInhRiszzs9L
34RWm6Ju3+6XN4V66j/Q3j6z9s/yEJdjCjzpdoXwBRm69lPX3MF55u1zfgQ7QELlGAKK4KB9/iqP
iTnEVhhKltP9tpO6KF3MS+6SpHYDqiL/a8HnJ3EVttI9nBGGPbAbtGFwuB7OEXN3UfwpGSZvDHT5
h56AM/NIwt0iXUWQmef11yle+Ldq38TmNIdJfDa9ZBTtVSoFt1nzv1RwWwnTh7YVp0u1QYyV2mCF
M67jj7yyY2EbsAZstDUmKpGeWpVUIdGe1C1J6GaSQQxvCwkVeuUbGhR3FhjbWs/AAqtGDUk2p8+G
KtcPZqOonFHg++ePxQDPc0y+/ObeGNCOp6blvUmyHG8CcflCPzB10lYL5Cxv6AihcgEPjebJuDQp
mPmFLWxdANu79inV3oBQi/uuFoRSOQn3UwyM7fgtn7fEBWHFvdMZrA/K6+TGQsKhX7B9OLKx2hDM
Z2THAwZYu/mJYYx//WNZHXZ04HjdQ6xHiWP86rE4B9mrpHXHFYAjGet6fjJL1Ehwk/Sqbe77rcai
ZNmbveWWCE4fFEFZAHGFpmcUnn2WFR5qR7rdzb8nbTHHQCpDXN6GRf7FBSTLoorpR5Wc7vbJP/YB
1VYxxIBMrzWFKnk6TYkTqhHSu9B+aMOYr2hjbiQDCETiMPTwZWiFtMqKmC0E9TXnamJh62vTMnS+
Ke3Q1PZCvVdwvJCXGZNmb5SaHV0W6UKhJgujbFCNjWxt65QzYiq6fIyrQRhCPPzc0q9+sTRrOfQa
b+Yjz60LtkTLGuFCLKRG3nNNxql+IbcxLNFGjIVEsCTtIEiIK9yULffu1+7Qd8qBLaHranEknxYn
bUFxPwY289apVAbXYp4AxMtuQHRl2Yqe0DCfkL6ULyPzRfTGL5MWXGvd50/aZwnZy1zbkX5R9A4M
wIOMlEdT6rKp3iYnp88P34VsHuz1ER+tsehKzOQeqY80gq9F3Aob3+AULEdI8WEqhKZkWZrUg/Mj
wguBoi5zw7PaNPEhmlgLkvf2P9iwVy8SR1XrJHBSyfrkSgHRiKNo+r+M2VZ0d+AUNOC7trdtDzI8
frvTfqm7Lpwzyk+6U+OaVf2RBNL/boWJd+bjosfoj3DXTWw+bprq/Ufqq9eZQC5GXEz7fNPCyfj6
BxB9X3VzPSYz990nG/GvJkSQRLkTgcoapAwbnDPdgjXLoWs3IlJ+yl1Ix+BN7pmHvnejdz4nC0z+
+QtiyHho+t8tBgbazUqi2+WdFXLL5yQ017F+euoSgtW85iQXvpDzdOV58O+2zVMGpPB7ltBghtE0
cM8/dTrU9yX+2sNj5xZwh9qrqEyJjyhZGNDne5fzNqpBy8Nfn7FwN7KvdyZUfpF+iA4jn3R5ANtn
pgXHhVl/d9iUlIZVs84YUm5PaEruZkwQj7kbAwj/iBFsr46QeQvsVxR4T/4WUiswz8BZNMxSEL6h
q+cZvJcYUhoQo/gQQxff+fslxL4F7WdoEhoA07HqN2ylEVj1Ki3RRvEJnbeeBoyIGiJ2x1DckPPs
zKxEeQCDkIO1rSAlPvamGLURfIHg4HovS3UsIIBRtjig6cSLzT7D+Fr05H8MXwuS7tUYHSfUrhRB
iy+GJLjYsQmb/4WgqtS3JZXlrSjPSp5Oswu7V6n2a2SsGX06uuHBVsdKNb6JOk3YDWRhgtPYbYlv
M/6Eyojtngn9MK15zSLj+FKTBTmrQG87YFGfEl0mMufrhlAzzjH8sQIjKrgj9Gr00wn/XvFN0zI/
PcJAt+njO4u83tOCfwbcknw42UKTv4b63TcEU3uAkyJmIWU2qq81qqOf5Kk3X8zsQNazbSn4tZPH
VnO9KGjMPMogRzFQiv797FqThSHdCHcL4uZQPUcr7Ga6JYYxpnbr86HPlu0F61PERnudtz3X6Y8N
V5oed4N0kZgoSy7XBsnzbYoNYJOS4sXm+6kGrvgcoaxHjsfZ0jliB7UEciyQs6aBTweWI9zH/h8l
gmrYfTtzVR0N/HMpA1NbOrufsI0s2oHWdCJm6bwuOtk2ug8zzbP/A39qJsIK+B6sB0e8qvEhjcKQ
pvdS6v/iQA38EJo3cPiFAdhdkwUoQCE51Sfj2jEMUjWFeVT4QaDqDxU8bgA2R9LpSHhqf/YSAAid
+w7iWDa7qzV9RV35fkPOJO1vPyM28AVIAQrvNkJVerdPyNZ2OrPw8hwXpEdYAvu9lKdlQmKotlaC
lAYPFS2nx6KeA8QuEcRM+xxGtLHgJ7xC4nbfNH1LiT9st00tCENRxfJAjPpd1Ukzo8XxYpTlBdrt
1112fcxXeWb/3lwzw5T2HFCF7RGUksG4X0DCa1VWUkdhY5U27+oe/cLPy2a0ftf9GWCvA6kmz+cQ
QzHOWUxVq89OFWrxY+z+3ZUxKAo6dMosgxD2uGLUPEMPnW/q5Z8P4KzWLcFj2ba431ZFo8CLCz3C
yUJrO6WsY3V0BhxdWtQNv2dpwgU4V9an0K1+92xAR0q1V/ZLuV18qzUYc5KMwoyAT9iTzcWYjZDR
Pr9vsam+sCWDZAWnXwqSK+3oaTn04zRj9jzE4oLKDeR1ZB8pHiXF8xX/TdeI60OsKHrrDMBYos1B
A+0tjVgSJ2ed8j1KwLp1tfZM0aSFNajL5JohgF6czm/IPYJEb6UKHgiOTcjIMz+fQUxY653i68Kj
lRsD8UM57ucCDOtFyhcUJza1/vniVKvKu+qyiw94GWf/ywFO3rqCfuGm1mO+RdAEeSuSaD0gvI/b
GdoWrPN8gwwtyo0+rs1z2RxAb+QdN58w9ZaLhioZ4S8+UZVPKeggwyNGcMvK3FZKJNoWI0tpAXNB
bZMPja74HCXtj9lSX/Mn8RwfgHqAceOycmmkY2eeqmo8/L3XM1H8UIE8YYEawUWDobEPfH9sluNw
9t9G0Tr/1EU0FbEZRCrNkKWKyaEesKWebB+EhDjdNXTd/iTq2UxMhBITufzW9c1pAr/SvAyD/1ov
FGUovtR0VJhM0f88UTJX75Ts6sxtl8nsUnZkwKKDW5nd5iFSFsUqBnjN3T+u1B2HWfzQAKVrjWaL
unD+vMi/5EtVYXAWZVz5QOL7/WFOOEUcN1GwmENcQo1I8gLvJn2Fhlo1B89WH4Ht3TegR1/Cbe43
G1/bv8r4Ur5DlvXOQZOkj2KqMUh0JovCXVavxP34n8BjwCjOpOf2LELlztSgC9N4yLpnh78wo6GH
+EmAWDnF7Y3/HmYzuL9N3ibgG5yzYVrQhRH90H75cwwmx+b5NQeMknkb7hcArfWHBXLVPzuR2u/l
tuCptf4XKMKl9YXA84hkqjtSDPC3TIXNnkWzrg/XTfafQpQMtcFllbPeMX4vJXvs7NDTVpYBSxoq
JpLWh5275cndGGaODE7fbZw/fckiON9QwplkVKiafq2lPZzMzpb5LqkeBMhWIO92EFwZrWgD7XPO
D2Dr71bKZ6VqS3jX9pVlx4vo5uRIz0jKeOOOQfRGkxBSScUKo0yhhc9yEK7uoso4En1QcwKHuNyB
iBcg9fPiCVXgmBVh/xldK56JRJyq1CVv3GPRASla8PvVpV2u1b55a0EPT6dSRsrhQXwO+XwKqOt/
PRC8lVPQ4GmUbDKvzhvrrk/C8M5Fhv0mvE0We2Xu3dpz88JfnvG/scF7IEkrmYxY0N1Ij7CQTfA5
1PG0ZMMV0MMtlvqJing1Azdb625Av6FsGEhdihz3D4lKV5isoaHTClylqtshL9SqSXQTgf3GvXtO
0+rWpKk45siFN52OhVrb/klUqbVAPdUKDiEVddrNRist24rNzLT2rioxQCyZ96RGXHpnj6x1Gdr+
Vc5wIkdKdx2LuC04lgAhM7pgGo2Od1U0gf15G6UHqEr/Ybnw/ve2G3SLuOmTUKnISkpItkvv62zb
qo2OD7UsPdeBsB4RF22fimcVvzLf1Kh3pOEqaER5mFXa0EUOf9zuepZDl7urGibP4MfsHnv88dXb
knzJngM7BYzM1Ynm+Z/fQIZJ+KHAnw0nnkjISYOvY8ROfiIOe2C1u/+u/2rhUhSUwB6CS+UN+AX8
qP77wzpAOUKQkwv3xAwzfslY7v6gjea9Nyy6aPasB9v2TZQmFpeeJW5zhARPSF+70LgRY0SnLgns
U1CRrCEuT7HD1kI8rYnyX74TdxBDJnVQc5R0qHCKzFx8csT3HeFDKb52AaDYhZu2txZqGw6ke8Ne
iJ5XbIMSuTOQCDFyZE/rCdn5fmE9gx5TmDGEd6PI0qpzqzf9A/5VV7IfGuFT7NAMZb/QpqBNVspO
yjzB3cF1Ut3vTUrtx3ff+2TVCEECG7+107dGdHTpwVzzFuabvq9ExzHtfy0D7NLeoV10IUTAsaIs
cie8eO2xOcHTxQOCIQGgaEpyVswP7Wvaf1hlMIVGQhz5ClY2WyKgnESt5G6iEj0g2dHahzvGGs/c
1kuBPrAa02BCQ6N6yQLWCKbumYUiWi3ocB0u/J5TzpaZH6woednf3r667I6j7QhgFp/ZaAe1hsL/
YwrLvxSHayMnQB49abPvGXEwEMt3isrbzQi0ufFTxG+4cJZVCBbl71BQZbQAMdTwW9EhqEoCC/LU
gDRcIh1JGtiNYJhYdkVJJMinPDLGATgNaowW6zxH3OCYSJ5HagtuPcRNC4XtgQaCfJUm3v2FJqvQ
hbSeIxpEolYFsok9rC3xIG9ULoPVbowuSjlN/tMCzvQZ+Ujr1+rM3YiSXD0btl2OA7u5w3zRnuhW
pGT7ksl2jSdWpAohU24M8D49wdX9/UpEG734vvNXyQ/yXH86JVMYb/olgXkvv6Q91GZx1Y7CekGr
tyaMcUk8UgGYen3T9YX/5fkPMNAuqFcDiHgAcnsJOn5W6S4O8B3cSfY43LhGshjD2QS8FiTRDObH
/OAJtFkoNjENw7TjjxYWyVI6IwClbyzi/azSw0W0GYg47A6BY5BIQJVepSpnE/7mXJFS3KzBPjqX
SQgaLrqtCcX4QLOWJ8ua5i6+yORR+ddhiwiCPK/keEoCozczOfpQbcpyjGFaBJ68Sa258HscXFah
pGuVR8NMWDDAQf0SV8sdaJvpov2dNH8YvhWiEEsVdBgRILIH3em+akW2b1JyxJ++R41DAIycb71F
X6FmtVIlM8jlbvVtEKUpjOII0WUI2uWwg7O5pm0LOxG558tSDewQMLZiz+Z7lMqGD6ve3Gekb+qV
xUngnxecStT4vimjzN+wpgojO3DJ+9Z4nF1IICKcihfjBdNdyTlGCd1a02MyoPlLh6JNrfev1XVA
5GuvftIkwct0BdwY/aV2YzNsM1/a7Be9iXASBgL+KvY9RsEwnuwg7jCJL6Q2zLG2ccWrsDa87IL/
F8iNZ9L92bYIw7UljBV9FLHxtR/D/4ZLrwerbXk/ADhqsoILw14LORc+7DgH24U4of0E8uEKHSXi
DfXDfcPBL1hZMLLSDrNDOoP//DjUm/QOfax6IoeXDwqpQ0BfgZxnDrk8jObbiRVdw28nRA5LL4zk
9GIU6zWJhXswa3UYhhgi4YY2QOo7KPMzYJhQLvWcRlXoAJM1sRKXjXff+6ghR3xA0KcZHjoUdelh
PVKNlK2Wc5dl8+bwrt/LRpXYmEtPMIrp1IKizDmhitqn11oU0K++W4xUZXkmHCB1R3FrKe5Ri+zQ
LS0kJf8KhiwkbjpcrgRokJh99eN2WTcNt0r0P+XJNqHoigX14zLN5TXTaX9xuMPb/uykWv1N0Eq4
fRbZ/MTe+5ZVee5yGbIu69FvrCFz2CeK/IBXwwlyPZh3KgroCWMvCTtHjcWridJrlgV+vX6ZS7Y0
a9qbcck0RUV4R9AIphZmEF4z68/4z09wk+TlQ2VPyGwXbAHIsW1UwQeA7f82/0ihkapzlLsxUUeh
eCP0YSP7NHbQp+QP6U2ybusL/8M5lytZqOBl9UkyK3JyrBqbKOU0t5CbEdeMaDikGWTVAPPSSMqe
lVClDK39xogH82sc/xr8XQtxxSZKpyJssawy0Q3yT9OvX6QrIc8/ChiYSvO1C5NP9NfpZlwaciLj
3LBWwot7CZQbAvT3Y8GuFA6ARpzy+z/4uX3FdSzJn2nUAYBlC4YPQVEiY0Zcp7WTflcq28tZwx03
FsFz41HdTq9TC4np5aw5BaPvT8M7joKQ4lDaMUV5muj53sMN3TCGcHppZnypP32723UJdFvD2Iy9
ZAq7k+1BqEfEN7onKkUA6/DvHsLvGez/TNRrwk6PWTB6820eS9JenwoOhyq0h6sNyMTo6GGhZD9A
ch9unoeDel2K8gQsP3QcLx1K4JZKposw896ZQkL4Qn3qBt/78QiY/ydc9xt8UU9ZT7KA9TPR5Ny6
ZDJh/1na7a6h9bgOe+t2cQMMf55pDDPirHMYly4U2SXZEW+QYN9A/8Cd4a2lx6BXaBgrQk/pPQkO
CmP7BuVEJG4Ljmhpp+Qq4Oat87Gz4jG7buc9j/6EHLiv13CVX/NVGR7E7G4P+X4y1ARTjFMGkj5+
oTN7HIQUWSgQ0Ue+MK4Vs2E7wpFTFTdzKp0TKC/XjX1KRWPqxLe0NbPRkiy/rs+uqPE2am7b/eej
sGkTqm6TM0sLpGHLNyFArkHHfuYiApE/5wd9JFkCBx/DX+V6lQ+D3B5ug1qfVRnIxXnAmEyWsBY1
J4Emn71Qy1lbK9fVkx13zZcDs8AAiLUO6BmB2+f4hgouQdqFcV9f9sT9HHWUSpbFwamZTW0aKTmw
IY5/v5nGFLs3KEUikvxiJoaX7jdb0ls6fCJ9uGTOvPI7TiRPSfMHamAtQ2BZLWXv9zN2HMy08tpK
CXHd7jdrMpVf84aneu3Gu5x5uZU7n7/UFyh1+kxQ6twSmS5gJ7Clp0LPZ6fH6N1gmcjkJ/kJw5AN
0AML98VPaqrC9pzhyvoFvyBnik2429vE6mKGlPEdBUgkOuSbbuEOGP99WZXsEiDm5T0g4Mue0Rd/
taGQnAE9+bA9BpyrcNDaF5Im3eRruE+pQchQK4KmTRVU6yn3YJ98m2ocuahvXO9nwbzRc+yHA5y/
f63OWXma2W8yrjLC5LRF7jIF2tx0EJhIJLrMPQZNSJZhJ5bLKPsChC09imXTurLRA1xUIIe1xbya
aPVkpeX5K7JHdqKXVKCgzoxo1WJJh++l/IumZxx8zsNKip+B7ymm4mPhc8ZO+odlwRbjo0eU6uvZ
qEZ0jwOpDAco6HZBsGYYhsTttYGek+iS6RGpDhgbWnacG+HAKonfcjbLKoxSu10EDnd8NypuIT80
jF3LZ0buJyTU7qzl48DRrF5MHP2zoTxYuYWWI2ZQK2riXXBboL2zgxeGZnbMYtgTSufF3o24spXs
2yBtf/TgoS3CDoAaaQ6LEgvndH2jP5YfuxdWK5mvWr0M5cXYbaqjEQYEAWuXOHl7nw5uchLr5Tt1
E90v0qRLyyPDeH1hoNlSAtulCjVUxDjJehF9PBagoY6/pv4dR23mYMYIDn89cqso75bXp/mr6KK2
oujhF2bAXLb/DAEjmcsX9IQPo7VNUxG5iOfFPxzp+5I9Dc97fg17vnXWJ/LN4GDnUoqtsH4Kk8xL
yThP5tSxsDYCA5F0VIrcWEGbrB9szlAdOoh0olyBBQQ7AwxwVTEjU0C4Mywu/6x7qIKhYdW95YW6
FqPBHkXvHDiAY738jE4goerx+mj1W+0A0gHgAFUQOsqMp1pYibOTi1w+VPqAJA40VYVRI17hiPQw
tVJPb0spXJ52c1gWl4WioPczWIGlVfDgSHVoadRikcyMo7vCTSZE9uz4X9wGUyIx3YBPT2tnF4UH
iBq67xT13tvztAUH5CPQqenDxuu442xpPTsxzhi1xEC+QTzePjRNihO5ZpWHHHHf7naxy44jc2Pm
VQK1kIFEOLSIGoh/dZomhzYWAOhYZOs3hemec2PX7uZBV89am6ePeloGMtWrvIoY7OmPuTNTfcWT
GtRh/NoFe0Z/qhrlSyNL30mPBR1ndVSpEARgSycl7wtdAF2Fj7ef8kwbZ0Bv8w2cjI0vxdyRdOnu
gX+MRUbiz/k1cLcAaDvbRqLL/l5+UknEBOEu0FegX2gnS0F7lhUQA+mmihcorod5NEPKpTqgQlB9
sD5mWFvG41LiLR/u1sldIn1UAfGvJtLjjmbX2eyOvf4W2O+ZV06deuBZx7H8gJ5Ct0EvfoBKJaZj
3+FMmEg3lnnhO0HKyMEQ47DU0VqAU6POIxVsHZF07Byh1myF7aUN1PbzpK5AbhJVEWhQX7E4U4/P
eGeHpwLI8nUUi4MzFtl474EXVtd0ytun24R0QMtBw9MHtcde31Yl8PiXdBMbmtVwBzsQMnIK+hn1
mgQXXehhYw6a6Z4An6ddR1pL0OVsJDjGLFn2RaMLoiEzQdbZqrsCtn4VBWfXMygGURK3zU9Yrouc
qsMlOjocYs9OGd/1veWT6gfKxQ+PSGdRZsaPGeAlApNZAbprUmyayK3OvU8BZT34qD3yTqphkA8F
vFySg8cnlm5/2h68Qr2HyXpJfnnqNWkbSDkFmvApqjHqLA2zPCvZQTwp8uc5a7Z56op4A8IdlYKu
oZD9glspPFrTVwUbc9w+utEGVHtot2mr72mrqvNtcYgN1YSyBQBgiCt26y/I5trOr2sefeTuIukX
IBI1I6K8x/giNAmrYbvqLbZmBERYLHjHJIvW6i1napjf9+t8UcCjcDMASRw9Qz5kCQZm0VghQMWH
p1PTgUJbjMCm83ncmnlONbZuszyOEgRN18p0A7dnnDeOAfsuSCwyqa2AVNDOKiSG0jkZgeSNvRxR
k3f0m1eLhfsuewpFkk7YT12SlW1Sy42UU+HzlW1xazH7QZWs+E2az+Rcsayl4EF079sb4EytNmux
DdwI0wkQ3QPJwaxZWg7Gg1IXSeX5uxhIUJkp9e5ofvJSvVTIS3hsAJQrRQa3/HroAWs17ozu6DpM
Bh8tjmwLH6CVp8nvO0yTQOSq/FDBImbqNboT5dXcDyv9jlTueSEnHOQTkL19XHJMlgqk0EmxBbKf
JmEwNCgVSi5Ac/f5XM16r/LEuFcfJDPGN5L32GTN6prn9WYYPs/e5Tsu/wfzVpIXjrOdSOSYgKjy
Jlcndn+RbhzGGb8KQlh76ZJQx1sgCnZOQiv7mAH4aqs/5IkTgVOqDyqXh/sGZetb9X1MABF89QRa
zoxdJX+/2iXFbNtMwMVtHl0rZGp97fzRvRAjsPOb9/XioOYBXX8KbHtx2DDidYsUHEH8bYbKPsV8
R/XHDs1EzNpc0aHNLw/S2wTJmDDDBJVOkRy3DSV8khxNfd4suoyTl/EXoHH53gi9TvK/nbeEu0LO
5tS7HhB4NZF0ZnQzWB5cS6eJhDvjd2VyHmWvwEzQHNgJJLzy2Qmv0LooYUcgcMTi1N7/Ipma9OtE
E1pQtTAmRSTD9w6edG23rQFwEJ6UeOagn8NzLwrafYqYcAPBuLUw3e9Hspl8Dus11wxgA6WsZOFo
KOR2BvZ0aLVWJaOVv4tYWJUjzMTnAKGSyaqs6JzO0OYZutoVVb4RTKGpGqQUZA+YvgBC/VDK9nWa
RGMr22ReSDOT1pIxNvY0vICUjx/a06JdDkroWZX65PkqbOhE/K/t1RRzWWQuwDVthajVCtdmrtZo
RH0jldKF8SMqwJABMdHKysR85yoH6VCSDYKJFeBdP/TmBGR//X8VER3p7wFVgIcOnvu+TsjycPyy
aG1TN3Hod8U02E6f+LGu1d3e9a2Ql8n0aBr2CFdv76xqGWc0vt33fm1F2dBHkzHfiKVMqWTt61dS
xSYnMwx4SZFY8umccoPEu/0pZr/g9AQSAsDgXHkuBQOkqfii4AXkxjKEuzkqgeQlTo6OdzmDv/ev
tKquKQNqbA7EMEGZGebVU15dt73gdzhFfE5CUeaQnP3yp2rUgYRunafdOos8a2Hd//KPOXpr5ugF
i+2N3jiV6YqNa0jGMtSfQecLz0z5AJxRE+T7UcRJgKuPL3fHqPa+BzVlOlgMvnIcXWHR5g5Gdka4
XhulpLgXnEm6WorgSZLVXdBtWF60CgRZ/ZbKB34miJwGZ/6VgeM4S4KMbNlG8XjvQI3gqNiHs3Yd
nWE2z5UDiFgPFDyzz5iKq5TxsEthSdx038Hu9S4IZEc34AC3C9aUgWmMqMoYY+nDnPj9xazMg1Ra
fUa0iZ+/ZPpuNx0owy/cazNp0mbaBVLVzsaNwPb68M3+vgj34t9FoVb2+MKRUYP+gkYTnuXapFJB
H1p4U7osf28EaHfcgaZjtYotXHA4jfIuoRRozUTo6Avr7Bpj8cEIWGf0cK9964GVxhHDsz13jk2I
OobQMxBUGBBH5/QUkcswMoIGS48uV7kpRyaf4jT0dtozKmclAPWyFgjT21r/IzOwRhyKSXSSSCM0
Dv8/RoqF+p3t/IJViAvNBcvdnFruUhYpbFSwAvnKGQ7qAuCxiubsIlQ9+8/bCpT6bDBcuIkQdBKl
Dso7Sz9Ee9T5UhdLIt0LllGrqWlf3S7XN4+o24So54HsC6Hv5uIdPLs565fUJ1dTKWBLHms4Xalb
aGzgzGWI2PxxvEc4smBJGW+c5Gy+tTK8SgUM+DRVt211tXUUUb48V5q4mVroDkLru7EyWlkPF9sk
E68h9n3qQnbhcvUhsz9QrX6pD6wk+yuI90yUAjb+ClnDbura2meSlNXu1YfbnIn/hGGvcwVS0uT+
uS+Wb/5Lyy6TYAdDdH7Vd9Tig8ljR7VC7E1YkRNGHeH8CqYCVEHfeuvOTGiVRaWP3LKjGetDEKET
xTr3tzXe/0u+sASp+7q+RbjaSC1zaLOWzBl403Hr7Fkn1nf5mfAAFcJixCGUYeAUvG4X+QCurE/S
uHfDdTDBQFNvvC+Q/Yx6G7d2mohV+97VJnCnQYn6v/Qb776swopeOlGKnmbi+eKmi2jiXcdZLLG5
kEHcgfW1T254/jpfK0AcJZYjVPm7IRT3abUWo+BtV5rqICR5gtLUHTiyaqGCZLb2QGw/HrxX+WzV
p1FIY0QwxKViJj5XN7NvmN5yOS6WCwVm0rb1D9JoFUq2Db8Truu3YgCDQHoEjqIL5yHjgRzta1LX
MChXAa6BZm4xAoZGbrRHd5jofOZl4rHphZjqN9flY70AJTQp/UPx9zrf98xkh8cyRimVxqNU9OZJ
IE6tWU5746zxUzICIP14UlrpJZR2f23aP+8xpIX2VbHVEK2GLb7IM5z7oW/tWvHGSxoQo8XBblGJ
1aIfyKZxk9S15VdrBANJdudDcFSQ6vtKwgASIN6Xz2gTx39V8GnDIdeerlnp3M4AZjNMwbz3CYqi
RwuRPTyFqkymkjFRHA0EQKhGyMMB1DZUoE/eIUnGQ4DK496yeHnAM0gW9fd+CKXGm2LU5iOeSNom
pSKREDSlNolonfWWNkCCsC0pjIaKUth3HZyAIpS+SjoehsCIFr8BRLqOj5wV1cfWeWlw4Nzn6DqI
hYU5DAQW5DgBVYKty+xkSs7UTft099J3x4zAeEHg1m6ylJI7GVpHZdtTyvs1y5X/DXfucE8v20F6
MZTgqpqL5OZjYDAk2REFTwc8BD7cYM2F5px/M5AWgCWh8FPjNyd5ko6qnlH6H/6gyMU8eKOm9tPK
xn5Cby+fSqlizXiH9E0gYQEyNBPnReR7BXvaS7HWSK4dpFFvljH9mLuJnkAylxSekQIrNDlN31/E
eL/2jU8AsZKIAuVSJXCpTipoOO/Ja1nk8VYp1Y08QMw91zA2sPBUHfRB0yMFszxRa/AeXmE4WTN9
ABx3x5cfzMjdp7Y2CLn+bpMczQpgWgs2avauFx3KgT0YhbaiA5zOTa0K7P/yADdhT2v4ladEd33O
Y2eUU6twLTi7PvE7210ATGqyHP3tWefalOLiFoLD/5r7pOgQBEQM+GRBR4hpbIA4iWv9h440Qgsx
mN5/0eeCG+7xoQ063GQ1ZcsMpufn2exGPOCpO2ZPmf9Q+TYPbGkAh6STLluERAHQ37k3VyxyCObl
JO42SUzpTRFVhD9uiRfHm2G0c0saamR2LIeG6d+qsW5hy/fpXhTTWcEKX269AVaumPzZn9W+M/Mo
P/bLlzx+JOS6QyQAMq3xGin0IS/hKyj6vfxgmDbgVKLls02kfE7irls8AzvnosZWmBhIZqdWGR4T
sDrRPrCovBB7+gywoAofIkGiKN4BQdtgsAsuX45TmH+uI17EaWVq3k2pX0DtQaL2ez15waXbpWMc
FBzDLDCCRXAmRmfIyRW1BhAfpnk55Dv3nT6aVpZbw702oUDjmei2KcaZlnwZENE9uGZzWDrKNkrO
Zem/AGk/G8oDashcPBzJPxMKdoHDcE3nNTzG3om0BWpM1OIdAkEdYEZWlaDGYS+qfPLKCwIU5jFD
RF4offZHMTks3cMWd4YgP+ctCEm41JdlR6+c7VZkPvSqmlhXkHJ6qCtJlYI72vGg86N0moy52THH
5vigx+iZP9KIGid/cAkzAZO27el8i83leqnSmgIN/nf4G2qAaKuLNQtQnmGxSUADKLtOisl5rDF6
/1bWTlf//fyHpBFPDdVv5RClOY1tc0YBQViLFleFppnTGr3WtzrY9I3ymbWOZ9bROCeSMJTHdVY6
VFvlCDlq+7wWzw3j8FQGVQLEVKIR6xZB6au6P2G/kv+XRbLB0I65aw0Z+cVcL8wDoLiG2W9Ozrm1
YwSrarRj2zJT6qX7eRvcojeuUH+RsWlHEevtL9ezL5OMP9yOI7eyuVdKB/Xfhs9xgaLtgP8slB9i
faAIZW51g8uT3bERzmRUkUX3GqUSj+P861DLHXLHC1xTDjNE4GgnAuwsx8ISlrN4XgbqHMJqYnLT
1SsDU8p8+yYFO5myTLyoIgJiCNy2j3gNqyKokoAsGX8Ssbic4LNZSnqySh5mxtGVwpKDy97ToAoB
pBBxmLK7zsiliECbkhpt1LY2UwiEEIziz5FRwuI5g87BGUG7KMd6J2jg0JclwcYUtT0eGtp66c6d
Z9Jf9yfcU7wrlvqbSMVn5W19Bs3gkh+l5mDzFtcsrej3BloLNGexEv5nFjEotxNFqXkZRT/q3iUC
jk6fZiPqNpdcVZRZFvw3ErnNjRhvR1qCHO9+ua0KXBK41jRhso6AhBxOfe52rLTYF3pqHbpjxls7
cbbKZeNbCRb3Q9dbjsU4V42R3MQD0Jjj0gvkQ0fV+mjJ7Y2OnFxC2IQTnsByullaBsT7DBeNT3y6
T4zTg/0IKrObzOe/aHqqWMfQAZz0LS2OY3K4E9WVBJv8hP/uwvxXB6Le++Suv5JKCbNJ5mt3ZCy6
jKQY2UG78x2mQk05h+XoH7qwc8aad8kzT9XZsRIlG0SDVLTdOWQxI4xM4udsgHY46abgf/IIoH9C
J5irruLP4dOpAuZy1q5lvcjaD6Cq8xb4XKaT6ARBntqhupXz18wjkNV9w+vJ/9ziNfzBcS58bVHV
BXgUOsh/OXzN9B0KBfzp7/C6vcMogrfNJJPBTkW4QxJjJ8i6/219AR3gO3lV7EEVjfOnirKV1lrS
Q4z2WVC2jiuD8AcpaDUGHrZNoe6L6J/eIQOZFJQfS18EMcsR+B2aRpeQV2vRYfuPrT9n7BOCaA0h
9tk6YhOMCfUQb3svUsLRezP92fDyG4czUQMMmGrqCTuW1Ect+viEJgsD6+5KZX1j86ApjybRsFMS
8XfF3YlAtF3rchfuVMc53L4eIl9LyJ80FSJ1nMeU4yt4LVDXT0DlKKJFSy4fWiqH7gOB6jLQO8ZH
oKxkr4EbLcfx1wtEZFaiY2dGDD4/kRFA73GcmbiuHo1owWIk4OnpaqL/Ku50iGF57nKaUhluQnMw
hImymc2imuyxWH0+HTZMtlfR6TtDsHPT/Hf5ALYq2c2bo6utHjOfnvsohV/XmP/S/qFEhNTe5t3e
NovRIRDNh32x18OWUp/7N+YkXSq+3G/TufwRK9ROKCdXZbPJdGcgiKEosK4w8vFqBHjokSAEQNkC
D1sc0RvyUYe6G9V7FjgvmWr3PqLCYX9n6QyzbbyPf5W2CqINf++um2vAlf+1DVP+GQhkCttOVraS
bNqwRqhHjjahagHkKGRSfUCsA1a56g5UeSWy1lTpUyt0McI51coaQxpdBeTfMHrOVvaNpC125Hfy
E67pLaAklbCvHIQTkzpTd+t5c93f4ZqxI92x1k6b6WPcu5TDqNSaetJazPEcf6PbBWaA4sUkwm0W
g2CGgLwa8ZLgt/FNFH5BiG1fqyEcwb5nG84aaQjsLXU1T8JrXZgTKmBS5NPTycrZXAx7fsYwiRg8
gEoXLM76q+qB0DSPj69NpCwPYG4LYYza9ZOYvKIVJPpFcNAfsUkwCoROxlufUJK/P+fOZUKzcWZA
zKJctuWZEoB5ypWAuoss0TS9nPjAyNFBrVD9GWxSitim6l7rd1tp8MDsf6zv5rhZ+hV+sBpckqAb
LhxJ3IfWqFrzm5907LkkjLUDKXKiiKWNSQnalljP1R8pLxniTVeqcPp1x+Sn75wCexShGiWYB3pR
7s02jHtzwg+DPr+SPZ9KCWZNLdc40Mi+erO1oojgOqV3mV7/1RTUYBfiQy5l8A4JxSblkGEIJLX9
oH0vOsG1r7dqbTY2KQ6qxhZtnXMcX1BTHojXeL+dDEhWt0RJxNKd8VKlKna42HEdb+Fqd+0UMEab
j6vbOs8j13zE0VgfxyMcYzmGre7HrDWIW/cyn1O5p4HAnXc6PH0OCXx/rxewBuahF+Q/AFjvL9iA
UuBnU5RVPIEtEfj05qnjAR8Fuz/WnskBZGKV39gPveIwzUI+zsRXT1Gqmknr1CnMYaftsmXR1a6T
M3MGX7WG21ym3V0Rf/8q+eoDxZCAR1TAkuEI6SAG/pQPzOC1tQdq9/2CLpNETz5Ert5BhwpXtvFg
0aoirt38V5ez4cKQQ6sOXnTvnmeBPOrtj7+9/t8oNMtRguWTRTkHSTUPw8Aw7GglYkNPeaiqbDCZ
pT7nKF94Ifhf8xfBCDAB2xRzXnfLHIYhU46N3HfKqu1etMxH0KfIgs2yJDGywxtehM4ZVrVnl5ip
vgiQ+QWp8rTMnurhZKLmumZfOw92uQXmZbBRDToHIJurzPebh3fbHuwE5F9hIdYgpWOfk7Or/ia1
N2O+0ICbiswSk1BDa1rRNFeZxhOKdKEdWCS3eY23yczopfWhkT8HlutCpva+aFMiAi8alfFA8fIZ
KujZysZp5yIw4LANpasTbUGtpQQyvGEIKL57rq3QtbZ2lAPwK2OJyS7J+Ek+zySsQXjXv9T3m0Jr
b58e5vV/KI7hBuZqRwTWRpCOXsCXOvG+++r80InR7dIa8JHFKStmnwyLTZVBIrXXaIQaJ2hCnoYi
HFWrbgGcN0hLaI4NOwx26VIRZ4HOFkRPqQBcV61jyV8IIc4PsIxWGM3uEgSgUn7aMShvdgDz6vJA
CeRsSNT/2o167Nn49yl+itwaShXxCLmV7a7lEJvnI1O1GohyWteMSCVb7k2kLOCjHGViwFgiaqk1
zy6d3i0mWoh8zM0vdvLJLhkgHiBh4C5JF43E+73tckPjwWMvH0BVrH8TtC5OXIDK5ZciDY4pQ4EF
bHDXGxML9Te4saf/yJ81/S3oPdvn8bV9jCs66mpY07mrNXVoTh2HlkZ1QVAmHkD8K/MhmCSutc+N
3721u8VaYU2mtATsAMGSwyp8iUZLi72VcIp3uuxhPVrIsL6lLBnqiAHuBG53lVfZ6hBvpNLEo0Ez
thTHqF530pi2va349wBsoZdhxLT1DCe0UUdJv9r+dvNJxiA8WenCL5VTvKQNJINNzdxz77MuX7nA
yYHGaHQfaADAI4fwHSki/1KThFfddJRQ4gVj+8xZFsQmb9tnsRR2dg7IMOdjXf2gKYkDZtXwkTtN
bG5Km/BblnDrv8djlHIRlQjTZiRdQvSxGjcbnQOeqw05f+CTgu54+ziWjVHfARm5b4xe598ssKsr
5KbSzpw+twwtiGsnSdWfbDoOQ/7clFotFnFYBJqe3ejCI3S8ZPi9DcTJj40TDaWzOxKdI8VJ+f+d
EiZguahTqZlLeM2dWX+M6hY+SIxyb48IvlB3tVAr7kSgROuDbJtw+UhMbHeqqDvD+DmQ+7GWhkoz
w1xGvDyFY9cGFx9QVR54Dfjv2N2rATPhb8ennfjJlLHye8G3ifKbRife01cCeiZLL1WgCa+BwTnv
LTyjPrhedZW5pHXS7YK+FNlw0heVcsrM9Bxvos6Xuq5SgkfSF4RhHJC6llO90lrLVwm9mZh6a2mK
zVIpq/veM2MErfcnKgBZiznkmzMgOVDnpMtPzvH5wDUwoMlHuespxRLICICuo6l6tcVfnMEanJrG
JaqlAyj9vEdUAu5tfQpb+jxCGV62263d9JD+7m5jChxx8molb4TSJ3qtZoFPUGmCCHWrMaCGl1P4
NUHXhcgkojlIgOVVI0hx0ghIBUgu4B9Ua2D34Jx1v4wIXPy0Vvjyp4AZ4cl9JifihqnVIwhQccPq
I7wBfuVCPFlZuVjnqwOICqc+rwidA5ZEm9CFXEu8gKi6s4zH3dOfJFcVOei+GTqJYd4aKdDWKju7
wdmcKAXtp1q9b3BgeI9cqfmIJaxMBvsR7MOKdkyVkguA2H1mFeoUrtVz4sLVJ//oPt30f13jYXft
lG8KMdq/00AC49EL81k5viAQEOZCmmi8rGU3nDWpFDHoUTJjuBg5rz7m9D49qCvZ7m+mZUfui720
WV1eTYjsGLOCb5ZQYz21tKl+RwiuMBo8BarKM9YH4yFrZnGyBMV4VrtRQXE1r4vD2deOcxtu3t6n
E7pCBzbM7M92O3m4sX4oXt8nhEZivT2va3T95sdnIEj7uaJmlM5KNZWMw9P3rnWkNbg+BIPusTA1
mFCHzD7luNT5uogdxowTtzmEl4iULApdGDH8ak1olzlfV7twtKg7KTw2n/7XzedmgywUJ8wep416
zgjI0MazhGUBwwvPb2Ckv7CtRCC8Uz/RMdUG/G4GottqNirgU50JopxBGswgJ8x72KGgmRlVwrfo
G5HUEGd4KUodBXFgMgE8j5VEePbIb7tvn9NJGm2WKPbNENNzIR0GPEd8H23ddrQ4c5fAmzht3YEO
IU2NGaLRAm9VgbIxKB1uqQVtqCWqEYAVitkUmpf0S2qZlByun8EIzJcLM23ArM/EGuzBHWsleEZa
HjG5DIkin4rM4Gsc/z1Gxjnt6d3UMcdctNxuFo+XSct4O5A6yHkiaBwVODuQ+np13hMC1rKO+qPJ
/VCjzYfKMvEFLX2VkhfP6fMYqnG738JoR8jUQEg9q8c3Rew+gvAjFq66PLGYtgthNe+KY1EblPUB
Zne0agwW9ctDCdjXy72T7sl4dAQLmWzzPrQeOirrYa/f33cHcXgiTeKqt12WLyK6cRIluXti2YPc
URmAwhgJhRucOYVx2pU/lpMTpBnjuAlJ7Q+sQzFQMzjoL5Bw5sIPC9EC+n6wWJeqeY5xBCwEuXxt
q9koVEaMxXyLDYzD6I8W4jueOm4xxx28eAllqIta/T7iIA7sIlt7Y+W6eOeEHlh2gwDqr2g5xfFO
KlqVZgfxX11ShxBj7cOPM4z2NJpgXjMkKC2VaTf9co8gKrF0CuLbue8tHh9pO8VMnjiuyNwsQYDS
pDpqa9a+HyZieMBb9EFfehCZan9VK6egn9pWOHm6ql1EaQj880u7yqfapMYm1RSOVd7VhmcHM9I6
u0uFg3atd2c2TNJ60Hem1EqzCBRWCaBoJWtar9wnPPD2qP2sWLa3o6xMGaiaMrQmmJy53jdRwmou
O0Q7LOpNSGNJ7Gir/8RG7kmJXb6kTnxo81iIjgnw8gSS3YhsAbEXNY/2sWUgYFu7KcLLzXjZQtBn
H8EweZETnKHoehk39reyhua+Fqk1BIWiMsgpQsFQ+AX/ippDykdDiU6zGRq5/D2W85+FUgj7oFcm
FPgn1v+7BdqNBZoXad5+pTZReJNH8Nx71lySVMdqtkA2fPvfRt5oW4feXyA+vl+i8oH8FHwNxohm
xIYnBWOz/VKNuovxpzIFwV9a4mllS8L4TN11cwiUqqclRHOkMCfjJy3kYU5ZWFwuK4l7SUO9oHTn
kMlYZ8BLUL5R3gFZZpcXIasB0kY4jOtC+XnVuCyLysR5oIdLfToaYwupa2yGjZTgnUsDDbJ4HrJ+
raH9+0v6dmp+ix38gWG+js5FaTeoz77gIdddhqdD+uJfNZum98vl53eROexWnoNsIM3fQG1k9YxL
sqRgrca5LSyaXUoOm9FhRAGe7u8wNFLJsn/WxtvxsVlkJ/jnvUZnkRxRaz86fU9qR3bkJDMix8uJ
n3XyMLxUb6AaFq6hhrxG3sXUiA07z3vLCO90FG9Du1ZbS/bTM1mGnFl/u3QfiTrexIblOWlKYmSe
hymBhTdctW2PeLYQW7cYV4r3zzyMirjzT88r5sEI85tKHFhg3gSadWmJlCaxIrVZ8u1rlTQf81HH
s2whxRvqg7JqF5rcNQ5jrEX0dxgaZm+tMfVH+CiOjDm6S7rTKfLv5/7I/VbBOrNSrQ2kCCTqV/54
TqOA0g9q3zCb0oJ8gwbuzTXwaHNccXEMEAza9njqwd29yoZkDBy69EZ/h/yA2SvmJ2mI6IHlP2UV
f4s+NXTVVpuLM18TAvhhjTYwMSb6f+uWQEyAKzn1jEtwGCmKYv9oq3YBb+8aTIJ3VY52hiecefJ7
hkW7PAtQ4IFCg4o7ksRzeVkolyulDRokA42Jm5Gl7K2oBlTSqvrLKZguApQuHh2OdFoXSaIvKQ8v
VVm3VFfZvn3mNpEgBGWglR7GxVxaebcbACzKMGlSOxA9J2a3kow18Dv8SA+eQsT8HvmvaAZFzjT4
KLRWyGm+22TkeAm5QxnMoSQI2n9Vyjgej+rPmttf0Iee6dSJgjrTDJHKKOOY3kv9cCdkq2MFfjKq
bEl8SeusW7uWD298EIiK2sMl22AhtQyE602b/u1zuvCWc78p4lQkr5YmavTaTbvbitT+pCQgu7Ac
CMKdtVm22zp/hWhp1NPSwldcQ1SB3+9I7NDAulpzo2gLUpvpqEIDHEaSzjTaKigR0O1O1anaVWCx
TRw73Ea96YtvfXqLzcfY8JWpBSmq+jHS15zPO8nd8dfmf8ltWufRJOYADYdWB80/kpQarGoQ0XMd
nnxP1561OWLicUjjJScxDmZune9dKNwH0VRwhHDhyuaCO3pY5/fqAIoab1OwL0B/ePomyA6GNlH/
z1EuRg5bMh1aChM22CPqqDXh8fsl8WaP5MTbQW38GS7REi67I3r3TwNOslRtuW2MkmWlPaH0PMp/
YmTQGD7XYUAPZJByvtNq7vj+6uRIyUJyVk43HS39TSI4aTX7l1Ru3rgF3vW6ge8BK1xPqVXmqL0N
3woP3u1SmQ220jaS6zyT/ErQQoVh8daM8yOEVh5ocIp4ADGOUBKgdlDHSC5TiAjD79RuILEL2JTg
ZgffVSAJKbp0+4yPLsuFrgEX9OtUVdnrX0+ewMZX5GTJ7vKHNdrou26HL6xCe90ufRwlPwu6s/Ci
lqXsIP1JMBS+jIGZxy/4jYQmSXsKBzV4+zbHK526XnRhtahEZVlAp1JIWfpdSp2w7wBJh7uUnNQI
DWWTLqxJRpP4QZrJgY2vkTLIQql9uROVe7xy4PEThKx0S61JgtelHNz/DpBTQRYf3WUHQ2PeJ0O1
Qb5CTTOhLAqpianSxdB1gbvjvPZfb+S72OtAatXzKkco7eTB9JqTmbX7VXPVlul6hSRHxDQB0jyq
YpB4rRY+g1gEg+nt/ERKB0PjT+RSvCGPGQ3ZwTP8dzWwdWVqkBgA2Y+fS0g/WKbLsTCqxJzEM5ED
zNWh6ADJy2NFNuZ6bsX21QdU51mAOWBdATADhBRsT9OqLZsBDwHKYxyj/E2ePgBvlSARC3dVXtsv
5ska7+OAjGVPX6FnMaTcoRuiNwV9egtgjep3VrFu+VrlGsS8VFX1Ev3a2TGwA+hFgTiNDHV1eMEe
0qkQZHX3cwlzH8lOh+B2CrzP1UQ3XKbEFJW1cHrq6005Lt9XnAXE8B9LDg0uSUCZZtibDGOhSQHG
MZYYfhHDfCiecfSgZX436FKsAEp5Hb7oHJ+pf66RwoSprSxUDc/N42NdrMu6uE+5HEL+rUJK0fzu
eLjMm6f2yPY3OCrme9xllsAgXUsKE4xsKRq9y96/zAu5NstOVaSEYVvQzN7FlznwP87VtqJR30v4
Tx9Yc+AHapGkD5use+3WGvMt+cb4KM8dDVt3KBHqqi8l3zqHEbJjSHKo0iSUxfC4MB0ls+rV2V0a
nzWG5wPU6us31sDIduAKrECLX0gOnEkPSy1z0E1k1f9dOA0wD9JEiWnRW5PghKphOYTchf6b5670
Zmue50FHKSYlSdHS47q/Fi22ratH3oxJc+3j/ZSqQ7ziDUnPQb2iC+L1mLaHWTXlLFVbrerPas1A
unrUmBMtKJelda5CR4EdorIijO9sjiuNnee5//RWsDAichyF0c+9CTu5OmjfbfwM5dWF1x1tWMc1
3zc0DvOhU+UGISlk5y6f5ClJOdFyXbLiFuAM/73OiQ9/248xpWYhWhXvXGwMRgA5YjIDaXOzMOhU
C1TWqoyrVp+gtB55howFkuiugJzQ5Ri7VgL99nY0BKrI2sInOCxlNBCKN0Hkl3zx5cpp/xlnN1sf
aEVVVVDTZzHcaWUgezsJqt+moHbNngX8kB8GG/6jj/DPctHa21FlK4lncN7bYCY3j+8P/etOOkaT
BdnWD5ceQsKBRwZIvMuQt45MY+75VFMKkjuwQiqiB5S0yMGpXXaQHJCrnc2qaCQsGoATSuJLZJrL
JAvtY9vcZCuAt+L/pz+yxLzelktrXIo/LiOPn/T5g/GYiVWbBYV9SBqlzdk+CGCvAIkiRxV0phzo
ullqC5j34bB7cvPhb3Y9auM3YWXCYGRkhgu8cMdq2PQneRuMFWTQmLxnF8/ykYePRYuIQ+JKY8KN
V71squ0oZZ+p/NlQlfNKcLQ9anzPz0QHhTEAG807vG7ta621Jzf9xkAb1TtjF173nAZd5K96jCuQ
8HvxCgOvcGiYiuR4Mzk1EdD5Kspa7Fb4e0yRDG+NMR9n2I6cmscGBZyhkW4xOjzWTiyTNstoJQYC
WM+rsqD0CYWic537IugWhI4pMRs2L3kJtn6+yjjJususALLINPpk4HmuJbYPqQvmx/TsnO4JObnr
H9/RYL7G60QQxlbGREfJgx39k1LCIXqVsxDyR/xVhhAL/WG4Tm0Os6Ec8mdfrBTzYQfqtTghaHet
T5opGHMcVNmUDk+XWc0l1gmDJxvTk/wJmttQjg/bnfGZOlhs+dxExOVt92ld88wEJTd/h/Tuo+a8
Ki4qeQ3IuhggrO4Fs9MJHBHimSSfdLx69FDQ1KwaF6RoWoDU5g0VYU8KJfIqxHWlP90lSZhpWvEL
uYly7pMo6JEVrEoEhcIKEzXv+Cw4cgahjWR+6GSTkd/RLmbRjAViZVRcU2XA9Eodra7E4ne7Ex8a
9Nkohp2SN6Q9gmOd98w7yCR4xRSmVtvIhB5cZLAu7V2Zw4IMvviF87l+9DDFF1qH/oce5zcVQ5dV
snbR28W/zQKJ30uji8azs1AicA09bBRGc46J+HgApuMTo1azIJsMOlejsvPC4Q3yy1uV+Mlg6K4k
HiLyFpowppmc1riWRKMBOv/g0FHtFNRYO2AvQ8P6pfjNQSsndZNfmCgOuPplRuEEk7JUjeBUd5z9
fYR1hxu5OcKY5qCilmFB9zHa0R9zM0nVypZ0pVtDlOIrnb8wR4i/TZRhzcIkKx7+H3kUNU4E7My+
7pTMeKMqhN8Lljs7H6KrMtMWUf1tooe1Wk03QFJx9C9jIj3DQ7Hgl6xks9vE4pdwGE+O/whvDsmt
u94vpRuVm/EIgiXSenWnkNq6BjMmBXx9t7Q2t2sMI+7dfx/10LciSYZNci1QbiYK5WkpWKvSPlJw
/aVV7DWFQ5dpdLPvmcJEqzqXJHO6PSY7y3I6oeXxyVodX6tuTbaoKHFy407WgKPpkV64oWN6e7VM
niHyIFFW7ObYzjV0OGn8G44Z8qZR+uAQ7h5Q8B+Yvgr9MqRvOVlTLYPSGqdw9umo04FJjlKa9jF3
fHBoPD3sU3qIMOJ6tL+0uICY9K2WrYHcb5048/rsoC99+1689NAXXtwVUBRNJvuepoEegalCN+VY
UTA9oFpY5li3qYDYOb7KPQth2raw1eu+IRNLgeC0Y+bV2H2DH3DMoH0C6nHrpHLAbR4LQWApcGGn
6WuaLrOR9esFRXXXSyS+75Eqp6/7C8LLQJT+ydpD4p5sewl4/pJTiPB/QW4zZ/yD1FmgmEGAr2wI
86KlP+6g3/as9ey/mz9cSmXJAEIDY0EnUMLK7k/ybYNJPROyk2A9Wn95Xg/hEPQ7uNEUDAtyp3yQ
P9ES91FqwcQpBd6NRhNX8JkFJXq2SzILJJPE7rwtZ+bkvSF2nvChhGvp3mDKgyRwnZ1qrFRPaiTZ
wvBnlGvR0UpIa2gVmeEpEJMmeJt1t1a6qP5NmgMKkCc4nw6+Cfj2mD0NJebP0EnPHRCqqg48Oj+M
A+2agexWRcOpWAelQP2OvfxSHkrFSFF6ob/SLlv8uzjqk6sDbaUVWuZTsZr1vI9CzdqScWfF1fa1
lnYitB4PakJU6GRfoZAxzG6WN0Z8rItnvxWzDNsPU6gOgFQvLY/oJiSHRbFdIRSvgWewsSyxTZqC
qYsptewBc9Wo1ISobkWLJhTF46mw4dkSZHPLU4D+iKxt2cE+BLr37j0759JFjJM2zOJB4+uUoVxg
VpokIYox2Yg8abMnQ5fN4zuGG56LlC4ufOOEnA2MZBRf/SYcsKyYFIU+humE1xQjdXEgoGBpBFRQ
MyJTDX8lq4npYvRPyGhQK3uRNgPxI0ReVwOybu8n+v04c4PrNdsW4w79Kgq1mQJQigBbJUjVtg9b
rApSVZqKcm/m4Z0+Cac8wech0bnQki6zjeBB67L3P/wRMDKY6uquiaUOFDB3yhoo137eYvazazVx
G3CLRn/nGtwwr6V/3e9klkhvYeUvFxp078l9blZt0e83UxmMqMf0Fvhmt1fGPWsXOJbmlI0zGWLD
XVChtwp4fVltO7tRLCphoG0M5kzI8Naauq2vb+MGMC5sTZ/wC+Tpr1X6Bkomaj5IsO3B/wW83s2Y
lN+IViXEUJh52+SqA5z37jtP6oH9pRydDhlPuoRDACZMZN5cs2eErtyphbGpYcZXUFc1kF9qyaMh
X+7oZNMDyFj/H84r3y+wET/GKcB4+3asVa09zzS535U30qk+/Xznbo/t4KdebridF/c2eE/x4oct
IKZWkCn/aQ9vkgsDWRgSJvHhDxjPgl9kN5A0aAGctZsqKbC6V4e/6RnzAby3f+1UW4DlxpTqX3Dc
CXP5gaVnt/tnzUrE4iPcLAqSqTVRtzLwyedj1C6EetgeD1P5LDUzJE0FoeduMhu7BTgDgYMlh/J7
aD64TZqyOqFanDiSgpE+nc/6jZFsH/OYh9YYnbBFiEZsKtGYdgBn6ZSI3nG6idGSBaIGJs8xbE0y
7Doedc0KZh0NfDQUycSPI5g+7dDQWbkEzZTi2spxOcl7cqAOXs8Snah+yAsMn1OufhXOCmcbF4PD
E3SqDZgT+7FjLPvm61lYm8HIRzUnC6+OKO9PnB8BEsYEl3rQLhRxfUVSfH/7YfmhHflWjUHouURr
dydvehxmfI6LAGuPTI1+YMRCL5eCB6xSddNr/k5B8lLCWdpQomBg2Hto0lW4FXcVMW1FWaRkUKvz
zdZyUDX9OK0TipcDHaImCtXxESkCd/1o02Mk30yc3Uu5MRcfaZzTF2/wBSwNCYqVx7T3F5hIOG9g
1xIwiCc+Xu5CY2PFHkika9JKQ7OVDY4oNpO6JQTl5J+EUBiFCR84wYuIQ0O49ilkdiPq548OJQdv
gvMrDzuw3mp5DhizPgbTaG6wMt+8kfPNPR1QVLC4QR3LO2JgB9SAqmGC0EVmst8BQERB6jOStB2o
u1v6FRSUqrRwFQ3mTIMJxPF2UXtcUdb7wACMN4FcmvBxY9TpJKbfa0dhJVbN+sjITiluSXSG3j3r
MO8t4EIDNFt5mB9k5lA4Sravoc3EsPRNfc6Ozvj2kx/0JmueEK8MSLX04VC29+nJUORNiTuR4nFE
sJnoziOkSBIwArqQIN+IAIQi10RJ9zYP+CMgyQ2/or/7UZ+FciIhXKFCWdvxmxd//dC1W5j/GvzA
YXHEPiHIK50EtPq8i8xgOvqnvxjWr5cWwd4+JFMcTx8JTYp9e1CgRsjY4XL/xIk1M3nIdt6m27W3
eLvt55nNEkkvJdSJrVTUBFjWCpFNSrgz+YYYSsvANOEBbV7A1fRIKRVOSoi3idPj1kxpIkNI68d0
mbFiHzsiwed237H+2Tdsl2I0nRUHb2LXA5Pt2XZr0ywZaZozpFPR703CJ7XjpKdrXDRdToYEtCzF
bnCrIybYKzGCrdqzHn4HQ5GGMAxVmQHsMf+dA/tgvzgjh53jXAkoYr6tEdQUwP4lhb14sUB493aw
sUzoczU5QtQYYVYqkP40Gj2cYhMAKF+7M1riw2kTDToPQff2k7EtJQLxbTk/UnTV4RlSW0NGNyDQ
Fs1I7PUWfzup9IAU+qZNalzXLeW+QlKWKPVfhkE6GnzK9qUzvAmD53w9jZAumM0hUtNeSzW8L3YV
9Ju1d49H0djcL/F/9C6Qwgex9VuWe4wzQWVXZJAfI9FtNGH2wSuHynybed8MvNE+h/dKJlsCCpmG
ScDvurDBoiw6Q/QhSOWyw5xD5UkPMtAzNByd51xHUzF/Y3e0Uq+5AHIaDTWtHOMpQofImkcva210
CmnuHuLIRrCQfspGL1zwrEEvINpg9QXaet5Ga19vzGqOq1Xm8uMCXIBtEwaN/3k6L306OQ2oimIt
A5YEGLfoHebM6L5jyGLDcCMKaxgTQOIIl59JVdUG7yA1dupwbRpr4Z8jKkJ0trN/ichDUvBRNiyf
TSvRS5g71r8h6HUkhLphvQC377n9+Q+pWhjukLwjxde9J1Jt5eXQl1KIkrwI3IpkmwcTzZNS5/Mp
EeeWLXFtHbYNN2rFZpVJ2f1vBz3kHl+xH3MGIulKVn3J/DPwkRW4DhXo7ZXPpExF6zGThNeBSlYr
D14rlgQhWnuwGftppRXaRXcG46/aX67KlbLPGmObXqvO5YxiRx0MMlE/4t7WtU5EedJ4Sia6gYM7
Z+Pw8j0prFqyzrKEWCQx2oskvfpbXN2HB01UroIs2FUPlAp9RAmdJgw5+4dl1k9L9VnoT5A2YZGL
3Uf9EEIGsebAK7NDbvu3dYXZqKMWQUKZ8p2PCwOQst//XCpjEO/8wXOLO9B8yXyvk2deG6BE/XgM
IlMP/+MR+uOr22gXRsRZADcmxdVcetE4Dwx9vBZt2Elc/iLXmBOs+1ZUfKqAA5Fn5vx+pSGNwSLt
QfbKujyA/Yz3OWDWVVJvzojmLFa/Me5WSPkJNEa38z+CAaSZcTAhSxTUTJZj5uJJp/3seIZjvjea
MRFumBV3QlP3n9dst35Pr/esYhg2dw3nqC2qsubtKpJb8fT3BMH+zhPns4+io60oTXEhhoVrULak
BwYmQsx8PeTcPSrnGTM/NRU+n70AhFb0GlCr8QbdeOYIEXEW8HQVrNccQIYodinMrfmPcPA3jfzc
8/HUt4S6PuSb2SxCoDm6pgVuvj/rHAWpcAvNLeQSKfyqi6bB8Fp1gDkh5nPbi/w0UoKCPUyJRmIR
2ZeDWdvn0vBPowWmP0uOmNCVB6eXw4F3QmQmz8GnxfrPZLoqZRVpFmVZwpjwwBkxJt5O948AdMe5
dW+wGdalbetpN4rj83B2RYu6z8uSRvp3NN5EbhMn3dyfz+tOraIsgrbtYIXBF2pzvySFYFqc4g1f
OIcF2JwmbKAFlBxnNy+AXTTPHChlWzxMsRJ6BER8zsYw0TCF4UdeWz8/F+MjReG8bdtkfFPtag3D
+FB20p3GYi+Vf3+YYKtQVtDJovx2t9gh4KbwdYCP67xAAQU/AII9s6YP0AoEx6dPLtYzVktDK9d/
eJibqaUOsg8XY71uMrJ/G8oU5bhlrRGqK21pbrZKvbLMr8TFp5h/cBw9PCCbxtSEv7k15UmNSaFL
jEKre5vuUD+ihJKyQFcYAkbKpWcGRA7Ib7dp0kEondbd7BxvWCuZ7tpqyoS+WJf+jWNgcXeDqHO9
4iuOM3pLfiuSIgjdRM9LuiPDLX5cFcCGTlOgN5eMDxMvXywUCwv3THtYTuaIRkMXBDK1wZnrRCOd
Fzis9A7CkWJnOsu7XEgy55nzgcnPLVp/pQHVHoCexomKFyt+f1E0ERqjk+bwGnyXVom+0df/UKUP
ZJXBOaGX4S6VdAs4IXFHuwRhCNw4DRz0uaZawF03adl6DHTNEF80MM46t1xbtHGLzExrBhaVQHBM
CkuRKbx0wD7LJkXtTUlNCDF+6vOA6vVjP7pIGCOCeT3ZWtlv8gbozOC8vNc4Fby+3bSPO9GPpv+j
EfR+IOGochfykQbXb0OV2nkBhJ6quScIy/4gfrkyeMpXYSpVbkzYuq3rfy6R0INltVoY6pYSUlMZ
5AZ3Z2IjeP/NAwz7qDUR69JgYmGyVk1S8ch45WDoZ5DwNrJfFob4KJtGkTmr6BjqrY9AH5ZDnhOU
PJjv/VoiaQE1R3+x8G7Cx9vQL2wGhENtzGBUYM5eGcixAnGVTlOoaxojW2xjfWtQ+0eKuKdh7M2X
HxLgbAgmFKVM22dDebBHUNBUnsrtmhFLphBSFK4AxW3WorAEtb4TxelKrMLTjtw20B+1EBthuDlI
M/p5MIR5Gmlo9nSxk9DlN7haRC8ChHyZ5uC8R7a90NvHLHktaGYRWvBYMSLDbODUg5yNsLzqMa0I
YEr8g4EbjokTUO6fC6VFlAOQLjBHohRsz/OBFbEFjtUaMaWQH68CzTTlTXUTPH2TN4ajGGiSPVRj
zY50vel5bzL9Ef7HyhQ79cNkmCh+vdBZs7hIKG/v2tUGMVOlLACy6K69E4/X8IseFjQObth4L2f8
aG5supSxciR5YsSzoKKU6VtgFJQ13Q8gFpwNwwunk9Cc/FCqRT/DKW0tjYW2iMFE78pkVv7M9qvn
CP7aAA3yXA7SQm/d3eOkFtHAL2yxaHzvE0DSMbChlY0mGiNKsMy/2UiYsQNdSCRU4vMiS1zjMQVV
UOKi0t/BlsqAGjP8K5ZnpM2dEdP45ZUKdigrbvivcVdRVfsXsIa4Ot00TNLPbW+OiF/m3cKBAwHA
oH1PItP3tzOnlsSgLbnZOhaiqQ+kglMtr3PjB6PUGFhYyfxfiI4aIaYwgd7eVXwmZPEH3CcX34Wz
GbqjZIMXGGMHU4wzWXpaHz3yxqsGHbzVxf8+nN0lS9VQlapfABS/mGdEOSNz2iUyJCn+ZrHoOZFO
+jwo6T4867jW0rER1gZ6EE5nP9eUvWfMxjONu/ZqLiEnCN6LxvxWB8m4S2UNKbPmF1ICkKcgDpOK
R/Q+CYPjspxUrw5J0zxySiRk045VR0XMvtXQBAukvt5trme4mc3Uh+evo/hEapDIEKA4RjrDWQgn
ShFc/vPxZh/t7iq4ZaqRhYj+PJaCnzefmsla4lcjL92wt9vdFXBo6+it36WL1J8ABq7TRbYZo/wA
u/KOpoFZVajvigX0JtA/UH0R/bPavz0lfpJBbrsj65n+ArRvhmvMtrTfZd1zAxvsxnr3pjQiiolA
DOw8eLqNd9g5A2ViF4S/noxc7vKKzK574umCvxz7wkkyWrsfVJV6PJXouAzqJVIzPD+E2lY1CPRp
w7DU5MO/WCiuQcq3uYvtyeESaHqH447yfkx3PSAR+2YbA6wyduFCq0uLQN8xPqzVOna3bFeFYdJy
WT4GxyjYuNb0eNsG7maHKklnG8LhiW143YNcGy1l6fnXn/nnHi1y5aCg0PyTZhC2GMwE++e9REL/
taweYcl907clAm2XehxQgDcWgMlTYi6Zk5y1ompcJjaJ+OVMcac+h8z7jja5cD8+3z6Vi3OG8otr
/iUTEEOY+0u8T6PYD1wNV4lvRzWApZTvhJJzmlpAZgWTudObiV5ljpq/VRpv/wZqM+bUQLP802I5
H60Z/ufQj3xWEULba8My0lyEUl25OlLmGwxBiTuDZqS5CwTsKIlOGMQmBljq5y7+1k3RZ3RWc7L2
OEUgP9713oki23mdnFNkD8+G3wIQfGGDno0HjBFem5px88/m0P9ule/EeTTUAlgs1QU7h6YTlm0x
0pX4c17feITkipAJaUq5U5H8Y9ZT/+pu6C6kmq/NBwgNAUKvDZDjR09yvbhpWg3xqYQPpcW83ZKC
qyaogxPwIrZuWAByMZyFVMZlB7XxnJv2dOWmUyrQgwf1cwqIyrEcsK964kb+hnFlM3rTMEmTuz4v
6cljBq130hgCD+IB3t9EdVLkmCFLe+DrRwaM7LCKiOYotlVq8VXd5Rol1tCgYoI5NlxD5sWRuMyq
vwvnSt9WoffVGgASbLcanan6crrcH9IqqcpYMi/1TK7isLAYq49nJK64quRvvAS9E/25BwntXvrG
O5ZeYwNx4q0fsMS1BHvnUh3RPprIYTCsSeci+8Jvjj4GUb61+/OKhHUR7KpSLWPfDUVD6DDXYUGp
rUZaajwh1RCbbkNS0qhdr/hpIvp+Hvbl7x6uB2RODvjdO58obfZFmONFQAFy2SoZW07LdwXhe96P
Kktg89bpSFgbs4kxyQvu6A9A4ZjHf/woVU+cQ+OY6F8eXbQymidbMj60NtJWIopFfodtNO4ucRlb
eVBsA5MpMxbI26r8Z3Af6DP8J4/rgCOoLr6/88YzJZ98Oeovy+em+PxGVEx2gB1/T6I5+th1ia/r
hZ9riEYuCJtnSSUZpvdCX0U9LMQHeiHbuZgfRALglJglNFRDokQep/DvitY4Bi5tjWHLyX+559JO
QqBSJZI6y9b7bpWmRH4DAUsS9eoYnzIuRg56K8yhwD8FctL5ctGm0oSGEL9X2cXjoXpbOqyhXI1Q
Y3AMwmlV8GU5hpdISWwoG4l5VkIaFi2qkwju/+tAzuz4rOHkUB0KYjdu8OTXAmt2+Eu5JI3MyQLu
HBZyTcTJiUrbjdysNuJYQRhimn5pd30Szwgm98IXp2BzOiApzle2bZ+wq8ul3v+BZWCzpRGpVH8X
RuTU1l6j4XA7N3QWIBGab+q+hEFAw0JInyoyg+UxyXxD5Crepb4kHBzSQsWrEoDbkF4zwETIljeo
z0qVvKxTV40vIPifOvHWYD1S6d/64BGZ9JCYUiiMr+4wd9MIl+L82IuX2z0CR5bf9gEjtIubIxe+
08xWvhZBCUGEXBt1b3DWxOQmjPYBQXryT20OYc4KdJ9WBa8Kmx8gYxHaxSjZ33Bye+tOsSLORM5H
CfHt3ETjElruUMt0sBEl/DNlIL79KKAS9cUzOPj/2p4VNPUPiTt2pqGeE78Z9+y32/Fo+pJdrGwL
ZwX76j8kEOS4h9A52o6K0AvMpJ2v6mkLODSgss/LtRZgijjXou1mjk8PpaC2CF9pj4IEjhjnE5KL
oRjw1Es/RgaTlYgIjpS8wco8me3uahnyKIBcRYKxtxK9TtSz/JzC5wLu1RwcbLRjDaNIHmm512MU
ljXHLl2gwDRwqBwnmmEdB/VFik13a7hC9s7CiO4O83VWQ2szs8bcs8zLeM9BiQlmOdI5j/mjY/jM
D5PakmPvfF96QCM8JWEonmQSpk8aY8rw4LpPt311TUumLBZpjvu7sACB38QMPnqc52fg4BeS728a
yXRYjV12FZhZpICM7NsHxwIJv99lPk41b7RP9EVBvXilafWLRSC0Bk5J5CLuz187a3QRaJkflugR
gCnT+fsb22ZpkGO2r3SqULRd1NdMm6vU6ioXXsJq1rCbVWBAwvI68qvaJP56+MeXMQkA8KQeDQXE
GQ0YOAoXwhF6yk6Ul+wWtiFXkm5zbxcJUpZFND0fDOVNNJwbH64P8wthqjrQ8pbEO+bRhtFdvtx/
PMSzl9Wo40tlvxSeoA7Hk+NAmVpqVa3PDckwvj0XJOwdoBEP9dDiJCpfmBDLA/C6sfbXSjBtaceD
zuARpGjenH28AUZW2Q/zX5mwcE72o10YJXe0cSFiJQ2kiL61B+vUGiO1QBNRokMgOXhSS4118GlJ
Y/7M7tBA+GinTcbZyuilXxjMQ5chdmL1vsdMlp0DfCbqpPtvx2RXSChUl/lnNqJQKxexVRQL/2al
dZNw3XfJxxmje9NX8zUhcoqJUsomDxTlIwSlRN9JgOLCxfV6c7Sn4Sq1ZD9Qyqac7v0vymb509SV
9evufImj4o+FBw2EOxue+eoDgmabhXyu7WWg6pa9wdQafJg2b9HwWmF5thqxuOIIN25jfMKPH6i2
bwiQ70/sCL/01iyGxLr/lhSuevIFjYEwXLBWK/1ZSn2R+3XUU5jv6mbLBokE7FM/OLQuLhSsjfAi
/CGyNorR8Vl4sJAto9d3566/8arBLjMhf3xWOIMMuQ/NfLhRxwb6kbnh9b48UYSFiKV0CfLIS6Xh
CGHjM1aS+QzMHTc2W5LvP35St+1F+b3fh1lNoysvDaUSJ0zi+89AfGzQp0UqYbMmax/KRMMALGwx
2+s0SSWzHpW+CKCQCnAbJbr2nh9emb47D78YiQQpqVKMy0bkwh+Qp7RVEtEYxxGFnQMhIMfOXmfB
h3LRJzQmOzbCtTqix3drHCWr1p9cUDE3wp6sCsIi64E7/65reeBGtnLprlt4uMNzwFRN/8k9PiGa
bDNZKz3+22ksDh8PyB4z0SznvULKSRDikXtKwKkNegRY3skPjC4WFRnSIO2mxwhYEp9IDbp++JZt
j6KHLZR5YhxqBkQdn64Bxjpad/AboWTcPV4U0Smcz6vqjI34SXTCPHn64G+gThy+GOfl3WWzP4D0
MWNhkOzKusZn8F7s9NavMOiUmYBywu2BErWMU2c09frGyYaOZZv0gwdNoeSI53FOP4NjloV5ecGs
IylzYTJFK+mkCV57rx9ZLa3qeboSW0ncPRy1j/r+mGdWqL/jR2WaZbrf4QfTlOlzygLuUBZig7G8
PUtLU6mTV7uZ5APLTNx0q5/ZkWwrSX5GOLm//empHnZYJJg+CNmPK+OrDGWWK3JmxTEE9aHoZDmN
LlhE/uDHL+ZTa8+TvOtCn2KwFh8k0RD4NO+7xxCHASwPvggbDohOQAeLIwAdRyA6n8B2NAUZGuzh
zd0AijbHbGSBobUD+Isv+oPgvNSpt8GTRkLfWTrI+waImnoQr99F79UwaGQxYVMzC2GDhD4bHA0Y
K8iXXhEO7tTtFp60O7a5Dxt/u3PCS7gRVJ+0t8Vch86sGIBilxqDxpsLCvSBBY14JdD/4+SbAC2+
vFLP2UH68nOwSw0zzWNvMa3KR3k2JZuas7x/NXLTBRziYULxrY94yMMLGRUDi595VL4+q1TrwB1a
Rn1PRFfH+vGw0WXpokruHcvQ2RmIufKhvbd3eq/UeRG11otbzg3I/0cuEPLVR/6rA8GtjfeJAMz+
zVrSaFk0f1DT1Q2ztdCO4tD31Vnxp5BteRxmIOtGZ7o3EoQScmuZQ+RDlibDesEPhoO9EmUY1nen
YcfBNDgBXXf0dbzdslA6X0F13lpo/n/hH0GArQPIBEji3o1JrCj2I/EFoMb5x8HdO/NMxq5LvdGK
IyNlEu0PMmucdmVXjOBOdHPMrkLJNSyKbE3r9JYzhf+UqTFcmkBWiNuPF/QDVn9OLFvUcORiYt2b
O1SLsQFsF2SlDtMZJAwTLnh3W+YsFu6nSbs25d7XA/f/938B4xCDKDTl7MCRNE0v7tk4Rt0JcR6p
vSvuRUEQB7EG8VSu6g1wdpAmdkmU4hbD9ngQgUR2WOUkJ+aUeXpgvkSa8FTkwEv25AQIYfWHihnr
v/DLAf4AOh0ioCUQovfq8cXBkilm9xrwWVJCPaxof1X7uAjxxYrLLv55VrBJ4tnedUQw4i4i3rbh
Q79axQwk1ORbPatNJDdYY8e7bvxDQALYGU32ALj/5HGlZk4ynZUdIot7Mz2GNLua20KwxE4dVePT
1rMG2L6CHN07XHXyR7EZRJvZbl+9Lq7fplKl/szlPwBEX/UWrsRAt1ugZxi0/6u0ji5IRSOInQfn
+EOZ/rsX5Z7PLU5N5Hm1/faRaszBuD0b0UCS18mjcQBvAA5DZXfVzs++Sg5AxxzroXxOFULIywSh
fcAPN9Cb1LhJFQjNQDsLsLuZWMaA6iCUym53aky/5AXmEmQz2W5lvJgHuDm2tny0e2iiszqwV/y5
2NP34s+3ZbLyJwWm5kO0NVtqWvuhEappURURaIXVzU4h34yO6zpO7eDdV7mSsLTjMCyHfVJsHpfP
wFaQJnKeGtqqy2j/TDKGnjDNRj3znj7lwJ/O7lhaGJJK8V8dOFYFbiFy0wSWH4Y+FMRncv7ec+M7
WHPnhlL4ZkdUvB9mOXqqH+1TnfkHSRaUbHe6l35Itn0Ym2tV05KaLYiMY90mINpyzHPHRZ9uewVS
i1fm4Lr/8fr+x6si+tH/Iah2s7xhEXpx0yW7pWli+bRYtN8RvEhtuMQVGq23O8rb15s8RJ4fGY9m
fr6y16D+UdtMZe39ge+waYylGDgMgZJrImojjkUbCsByEALH3lxkQhsasEzv7HeR0cssQNG660bK
BufWM2/T6/RFmadqCwjvptvmcb0ABGqksi4ZOGwjRKp9K09Ne0F0wDylfzAMIw/inblSKSlwSG8m
lDwnecJWYF4q9wcYnV/yV96wqwlw1K0vNAnpQ5ENb8u/OXFVjCKZ9X5ZEmneQ9IMBI80ZJam/m+p
RcCMYLY7sihU5GTj9A9TOd9Rl73pXLZmQe2r7+Th4Mcu3sXRzM8OnGfAhOVr+o25JXWsRvtkLEXl
pOXBycT90nLdCKC04NcVSW1nw5bgWX7zPsnehNiKlipZ1nXEooSma5+iBprundYVXTRIRE0ExSrK
KITaszZsRwQtXPnjJl8pC35RobniUVlQ2/noD7zafuICUPkgEXIKsyD9qsuSMjVPOEGs3v3G7JSm
y/n7HWSfzVNO8vjMtbQiIM/ZliBGiDG8a/Lgzoqt8x9c+O6+Q7E099q5mS5QtLvgki3u5/ajsBAu
G/5rz5zGxFvgcJO7/S/uGe8ynoQUBw1hzS/3eCdkTbqbbkmSG4aW6oTULT/v6bERgukori8NldS8
lXSxgZZ/J69AOf2tNs6nJSE9zWrkNmN+QXokJhZoUZRLg4mLb4SGaYiBgoNWpR+HkTsOarciUpl7
HcFtYPtjWXNAb5rjE0At5MF0ztclgGffY08k32RNjzangLqPBNsD1MNycYY+rVtU4GDjB2Mo527U
YogzueJ/dQFkkvz8ma6zNi4ChNv3Uk86aR8OvnFuGpIzRzC4TSMtyZgLuhVAgIaK3AJzNXQlRmMx
K1Sq5+wmYcW5w3B3eyyo9gju3hBQ2jtkDouSA0c0FogeezhsjCIPvLq1b8/BBXT3F0S5TWdn3Fpw
1I+fhC6lZpN/ncvVUva8a04aPcdmfJjAF9BIazpujF4Wyma20pK/UjDMwZYABTxiaU9fsfe1GaVO
AKQEAB7D67exJwebD/rZTG+TYhG8hN/adhVjKCEzCXhFNq6VgpAoX4YYy9hePTI4D4yFSkxN2a1g
IHk1n63wiUloskhzJi6HM8S8XJAjZfTFTbd6DJVlz056Tj5YKOx6nILG+cbsfu/uwZw1D00BVjEP
qbExuMOrFY4F2s68ZV7nCrGE+eouvgLVVDxVqK7NrXs3I7ccJoIZmxrJ6Mm4cQz5fCKgc8hoM6AF
LYAxNpdffaEEQaZmGOdRvCGLAReQ1Q/LHB19CBFfygxl6T29bSUJua9ASuFMByFrLm6FIKFKSqa+
h66ydnOIvIc2a9SV0+UxbdfmRZkmhFcq6vPFmKAcIFHKL1GFqxazNdzSQ0rClbDo84enRCUVRa88
n0s6BdEeM6K7HMLv4IORyHM7iKSMw5FM8X5ByLVHlSb7wctgtFVJ1RffCc8rMVmi2on3rWql2kJY
eozQRZo9zstCcdldvSjRtxxTIArQiigqKwpqEkIr2j7OzZjImRqURn2o73V7yCBIjRi7hCcCs2d/
+dG5pQYUQyn5qZ2Wmw7TplmsSJpi61LOluQrdRo0Z5HtkmBEO8DFcTc4VmfDbuzY46ruLWQdRMQv
YGsWMZU6AhOX/uI+TXaJhkDGsg2PUsbk6iHFAv6oLCflHS/6N7JB90UrYCubmrMfMmiOZ8U91pNL
uxPJkqG4O1S7SBbdBSC7NmVPPxvTG0Q8dJPLkoCWbzEBsAJvnxq4ZdgzuL790DLAhHWpjP7pX+H5
Ntx9J+Rg/5ZH7196a2u5rrLUvlC32MMO+7xXGhGgOpZvmWZCX+ADuVipryD8A+T0+vqJNqlsZdA+
2bGkwOOHZ6Cqm8zjsEUGk+XxiAoIj50KFHWrO5ANXqwVqFS5Qos+3XtVUzkt65Lmy+y6dnBpGvEy
f45wNiww9/c/WgTuB/JpunGDVm5NXb2MpJYwY3V5OniuHxB81RulcdfNPgzhbo7P6bsnjZQpKoPz
ylS9w9xepKVA+tVGV27LcpFR5CLiUyXxrlU1dIR+Oz/hvZ5hEs4BQ5uOCGioPvFIDpZbzXELRBZ6
TUNnUNE94ReAqVJkfm/lVMXcyyExTktzOdnNE+4Cpbhfzsee7wnc6UD3aDr/Z6VrSxAmd2hFYrMN
vaQITxHPWs9vYf1Eh1VZaZvu/kznb5UcS8Yzs9Yuz8r8QHWhJiy+cHgdgmdb3EnPxs0GSZ+c/Fvg
fVCXt2jm71yii2DQx7dv/VNC4a5VupyOaZnHjQpgvELQUtZYR3ovA+1yyzq1g7W2AxeEQT5wpK15
4wztwRF0WtnSVg3VCHByrQTPu3enOHtl0HIIR3LaKxkw44D+3LBqYeq52+7fjfUmWsQB+uoLq1sk
bHmTNzpXx8abz5VI8RQ6MKVP0JUdAIzbB+gP21f12vqZjkXR54tA9eUDdjNO+f/rfSa6JT/NFlVd
uGMcgwaHQDBdfh7RGXN7/t99H83QjPow8M9/iPSJUZ48N0OL5m5J8DJl4bEpfE66gNpkpTy95FUu
Cb669ye04VUTwCpV7qINDSyqAz3rTlsKlM7Kdtl+Zq3lPzq3ybKYo+p0BArOJBod07qieh5tEW0C
U9t5dWwWaR3mfiaGU4kGlJmFp2T67QlsAFmN9y02p7ZoQiOCsoSzyk8U8emKTeaarBhu31VO2lxF
3H4Jw1qbcyg4c3CiVGEh2iGr9oiIcY7IJElMJQPPBuZVTBjO60PUXfU8Gbm88yrLMlFSgmE7JFDL
gpN0eNiXcDEQoCgJ6DNpiDRb/aGY6qu+o6V36b5q+82pDakKfSFuX9bxf1dp90OB2BNf+5zKnQmh
08suBKid8aYgGqgW7wemu1vprwrzUXSWUr53lBoyoDMsIb8Er8o+lbI4jBPQRNSEyHblxwL31zHY
F0sycDGvzk3ox7sLIznHHRO17olumVpn7zlnOM6TVk9wcZCQ39sGipYpFQrEbDD9z++1qjR02EzX
f8yPnMITy/oLr3jGyXLO9NaOlSRnDKlIawgcD62Z3JP2zCcPAICZ6hAM0ZS7mYK7BrOUG9eTNc1D
S2NOY+qZn7R1/IOBWhZ/BGDfiUac84DfXJreTm5EbknMG0/Gv0d6JuS8BbuKoP6HyU3plnGZvp0N
6la6i+dn5fJ0N73cXM2gWF+KKVWGvwAgBZm15ynYn9yXABV+iqWwLGvzQqe/ON3+IhQpb1HxiYot
c/giIJuuMnbcrZjow4PUdyVfyfDwOhaZMFuNM266R+8lnAJvDqPseODx3r/BUm+4CPRqBQY9hTzt
nxmPgZBjhUmENwVwW6NI7VZetcuxkZu0iGphYtOtHtPnF6FYsYGvh56Id/hR2rOJUirRQIC9PzY6
3zhqlVu+6lvtT+yODiGwtTET36JlKOXhXyx5VAQlUXY3MfDW8AVa07PO6If4V3Z0lHvhWhG3B6AX
Pe+WmoF+CllCt0+YZg+ikFVYUmjEyTSuz+r+5oudV+SXLJpK+6uMdLj68lFvbUYE2icsYSK/Om47
duggiuSew4Whm9rmrWYPqWqnAycC0RUOyU7Q9AlG5FBKResuzti7YK+MIcjEKPNqblK3HXUlEBSO
VFTsi6ZeU04x5ByhVr+4Nfp1efcu8UzE7U30TOTFEuFygMOHeQHHU17uAC6sVpy5WWQvtBYDzVEZ
BbGgXRaqaMnLxhfPjtlxdqXrJnBzB/cxe2mhKcYFWWR9t3IB5RFXpK5bvhOK62P9fjDhY+JUZC6E
wJwr8Z9mA0g/ZRoKHvVRqRHBm2T8rNuCY8/ycXJqa2GMAp8YhEdCL+vW04RjGjWzSE50E9Yfix3N
+jI27CuvnlKeqHTfuxKXSKt0EhBkI060nE4tEHBqBBsVa2LGOueLjMrs8o6HeVumj7F4aMaY0x4P
GpVDtyoCSQej76uk6BylIg3A4PIMMVy1Qaax92cq1zL+RMIz6rGJ+yfSWY4tIuLaNhNQiOCy1XNI
Nq6HJr8IbFFq+MiQeCt6oJlSs/TtggZd2B1jbkKzHF9NajeK7ckeYLLT+O9sXCq5GxFl9GeFnNGd
VuitUwNoR5RzVTHOZm1gCOBUDvwVpQxd5c1M5a4HhfU91agl7kIeBr/oN0rkRq5s/upQYN5g6IKA
evlwc0fmSo3ZTd4tPN5EwJBKBy7dAYrVCQ8p9MtWfzpnJk+iSsIpPYigO9BFatXD9vp19uO1RiQJ
JLON51U1QkdjeeSYT+XbprRHGbaaL5E00+DqU61n3PQottw50/ByL5iGvL14bLFBgnrBbzTuIye3
XlAEQaIewEUCL/noj4UZaxExboYXQU3uRcXxGsJ3Vh2LV1+n+UMW2l8cOsjJ4bC0fRmrQ3/eTFx9
mf8Nw1Qe4va3+KHkztN7GGX7z2vTj+mnP3lxrlkFXGMa8i0gkbTnWvKS3NXA74plytW8utMSv56B
N4f+DxERgoG4jS1BPbW0fIF0ROBzDAyEubZn56/N11hu67YogjzEjg05VWEMQXx+HNyF62bVpNM7
jejIl8KgvhKf9ijiH6Ru5EJ76fNqn5QD6/F1AlvNH8gPr5lunSWcrF6I7HQvCqe3W3kS2h37KP9L
5eEa0qzPxfXYn3bTZOYZA2B2Y6NipiE7ZChW7rcSvde1W7znZ37A6t9ne2C8DqqBjdaeNt0dO3g1
DjFo8rEMCTUOJsotV98WfeC29CF8u9pWUYNI5fJF65Kd9/+4DboElXbmttuhPzOm8ECIcAvULvwD
vWF0VRIneyTFwu7t/FOCo9dq1poiIiborrtotXvBUnxl/q8nqORe0tROhBQG7xO2xAz+H9ARGF/1
qlNYqEaibV0pOSD/nmPOcOnrBfMDXYcJY8hqJ9LH/j5dclst464P8Hb96JMANXqEVtA/LMD2Dc24
pFQfNpDjsyPposjhLnqOoqXX2VvU24/RWJQMfTr3I2oXxZ5omNhxSTCtaP3Wz1j+CJqaY76al4M6
d3uitRs0Cty0JjXMz3iumu1/kqN/JQcNm1E3EaOfHUBTxPPJ38qyFVTNPA6UKcqwqh1Py1PsgGD0
kqXdzAh0PTqO85fxYhmpEpdtyDw/ziWxaRyy98dbGgOAYQbCeEQw8VffCmz2xplzIWps5yv72uxh
EqR2uoZEz0knO15WMKNGY1iBrhmdoN2KnOub5vrV3Uf+E/HdUfL82l/Vu15u46hqSnPlPk/Jm7O4
H8JrcRnH0OAjoZnWfhRPftnh3hxevbKsPaS5p7ODDw3oXPBaV2mu4INtZMjDgC49Voxbm+f9lGHC
yDTVXnmrK+3GyKyXmXKen8JTl8U9WPMWxBs5k5Cn8a1BNr6wRT9o3pI3hztgp8+DzQMUvvY8yzls
X4BZl6zxBrwUdiY4p9efEn1Y8Zzb6/BsTaTBDRqlJiPz6jxMpKzFEwkYgkrOAT3gDma4DRRge5p9
4lm9knXrs28rtzovNoQHrNi165hD7s0G1Z0ms6YZb25P6V5Rdx9FGMNhS9bt+e4ek/SLZuGR//tq
uAh9+7u5WotLZhYtSJ+AtJF8+EmIgRQUFHBDK0WbZbUwyd1osGUbSueqUoJjdUZD31Vmh1L/ufg9
5KTAgMAo9Rmi1ezRdXc3S6yaM6gjaFzRGzHcqycEA9qxG2uabkO8R3PMFY3Efw8hH72Q9rg30+Ky
2cqE7oFT7u3K7+JI+H8JCJnclqsEM9lDPi213rsJBmzUXFSCBMrQeMO7+K0PC8vr9lW9M5xIj9vg
APthjsP2PXSGMU2j6QCIEVcUT4eAl15Yp8jHHjjtDfe/MkhYMeVccRAHRN2WFHCiuvLu4Fp1e/gh
h8fzWYkbLdQ40pS0wyjVKcZaJjz4vuVB9+ITF9dFD6lf6o0HdaSOpSyWQ5Qxw71SUYc/dkEnGErD
UN7OPDC7HWpKVfPbDin2V6nc6R0X8xi1Iv3/Bp4mHQBDLFrAVojEU+tP1TzCimeA7qYulNTxMqx5
32BQHAs/S1xKQEOhOOgHN55s/Ku8L5xNS+bEtrDXjtt7nng0tVhXAkzGsZoHZZZaC0FTOsP66KfB
1TeZe67qDA/IekD12lDfJMYTO0FkRtwEeLAIZr+++bO9D8Symg+nniRUPVvm4wXn2c2Dpb604VUP
dw4xZf0Y4izVHLIypimlf8sFow4MKa/YMVEzvSmUpZ6zDQEASdXKFBgApGI4QdgZXU1kMgw8C3C/
lqvZlzjnIT2WqilDuM1D7C63j/7kLHMQhAxyhG17QAQVq0DJ+6HM5q37Bml0jlrXPycJCS7UJuDo
UbfgIB10kzK4ujeo+f1cR+OG+QIfSQhV/KRRtdze16p+OSPE529qgS5+8hF1/fpdlkpUL9BeHBFe
n07cTYSXUeOCZZ+OXIn8uuPMP+1vk/mP7FV3qCLnLorUusZR4b1B/UHxcSc7JIayuYfzFW+SRpDS
fJ0ttztlWuEvoYZqNYp0HZGA1tuXCpolaBwKKCbY60UE8J37ER4wyzaKHHM78hz/wNJtb2HjyR8c
lo8emQl7EgzMD+7z0jsPTP+us5uDvadqTCT39AFFTNW3E4e4DTGRPhaURYgGRY8yGUvosomFc0ad
gibVFyxwLPtZ8KhKS4vy1j/7ad4Td7g1pG/NHPLDsuAmU+ZuphhF1Hlfp/sRjNq0xhv/hsOiLlre
GQgfR6rVd9gpKto2y+VkGX1Yu7u/n2cjB4OKoG7gIgpcXfV50Z5q+2wu+VFlHGqP2JoEnO96pvYq
FALWDxxb/OXBuZ3ymMGkpEODXE9L3v87Mt6yrFluwiGMXNIusmB5r5qY4w/nmqfPQ6QmreYbcOMB
OPPsAgAOHAX9rLXW7H0czv+o1WzC3qvLNtiG1SaJBfUhMzdF7jtCQLj2BwdeTF6eWj7sCJZ1ZjCU
YItth279bP15vMRVWz5hogBcpK1tyZOyCEeKQo6Ki7tyKBy66v4HC5NTLC2zEgrElpgVXBNLvVDD
iug1PB6ZXjPdYgzj9bKBr9hdCLvSWR+KhJwIYsmkUnvMW9NzZV0fZKQwwIIF6V5oM0VKEkoVSwPU
6tZsE53NcUDZdXlYun3Z78oQFdgS7553EnMoF6f6hOxDhJ3r18vwX8eVmK2IolkxqBWxlLKd/kWC
zkY1NKnzMbxiHTHbih3ud4rJKrjKFIo2pkTftVbknGyX2Tg2h8SaL6SPCR4nM4UOHSkz/LXZ/uxm
MA52QVCA631IM43VUr/5qSDHmKBUqYdc7V4vHBUfe7OJOpBUjinauOQE0d2zjVjTrmBAQu6AMUJT
XfbMn0lOtA+7acDzPn707gAfqOotje+zws3xzfDS5IKldpOBi6COXUFH+DPLvAIlEfYZLReQNsTo
poOLUcyxHnZiu3xjGjE/VVxPMlzL6Yqb2zUsB7DIIkEwBkcW6OrAO1mOv41qguvFwyMK0t7JlUWP
VmYxWSnT84E6Vy8X1nAn5ZI1k3udhkQLZGPmIjqOHmyFGHVYBzYLkn/vkd64uqpoClY+hiFt7Zoo
qjBCKeni6xld3Luh7++il/rrSHa5R2474IQX7ih6S0iSM8SG6oMujxZrAn3j8ZlQu8V6RHBrU6W3
8x0xM3W98iV0/4Md3J0XDKoBSfmUP7OeDbr/hnm7zc8AjTPRqoWq6Vfbeuw+iDygEKtLT1jfJtVb
JTtgvlUfTKzxTQgfuhHi5JHuBECtFPyM0tzJGUUHMk1RDt2fygpVdprB0LxzqV6sRTbW+Ckoc8+U
kGQ88kIorx4uQWDSKN/qN8rXWT3Jdzbd2nVGlkPQK2oXIv5Oqu2p5ci+ueLosDUDokq1ZJDh1TZN
/aW4xfACaqUJxxFQ12BdLGcyymX0NXDoHJpqvunQzexNDsMRJd9XEz97JUII3CyDzC8MyuNdfU8Q
TVFwnX5GtzJy8FrNlJnmLAhOdduIobPBBbFmseRU7kVQ2OSEjZTBsdCJgcvE1IbGaG/E8qQ3/bmn
tCNuYXH9knO725OEm22xUm0yn/Sa9IYnzIXiOglndPYVOfSo86yacKCni4VGIwZpNVouwW+JRA7C
VIPgDtiqLoj2SAhQRqzWJKs+W9Q5iRzXMU333O0fzdxA4AKfnNpmK4kzCRBTNhIovcZPQIGl30Hr
1bQr1D2ncVsksEZVOAjm+F23ooiKI2tYqeMfZ5etJpvqS1uxDKBGpUd0CFTWo7S69oFIc/lKCEpu
eiOpFvItUV9nEv5C1dnucmxTl3tMlk+Kst3Zp1ayIQqxcTdNa1bZ19wIWIeoLszifIUSrtVug55/
J68KPb00X+UXgmIf3jcqr3wv/o4t4nznOzqhrbh0rWFUBDhU31qg86TswTROrSfkkx/rjgWGgvSL
Z+8hjNWkRMNQ/OUx5moXctaVSJ8R70/a6UC5/+9gMIZiQNiys9AgFIPNl2Om5TIn03C5Ve+p26a2
6RBIyo1n8yuLyUhDp7RGUsan7XPF+p6npAdIJ4coEeeiqD0A9UdnrAy3xn7/27oE8R+htCsQ31Sl
Wb47gi8KYlhwZT0VHCmmuBONf9ZdLrwTg9jQMS5VPxTf1SHb0O5hO63XTTn0Qgp9nUrIcEtiP9Na
kyoY7SV5sPOnuX0FCpYm+FsMOWimgfY9EE5zfH7Fz74bRULKqkU9HXmDvgXl8r36xaVXkP0GtMu/
yUe6i5KUwOUtEC7medfn6rExXXCjbcYgDQkF6nXpMxmxus/nfyKGHQ6fpLnm6YquSpQzGTUcOf0O
hm5+jG8sZUj5YjHQvX/zZlCUoGb1e6Y6q1HhfAysMjQNAg4E8SnHo3drA/jhQ4ytvMROb/DUXdDp
hRciLLJQWsp8E9rBfuwRUoZAyzIv/ihw6KZYL7m8MvoN4cdUcue1ksDBosV7UjjHEu5wahez5WWB
g6893epx9k4hBrWuN+ZIMmw1dvk4rkeztK66E/AvjUPtUB96stSRg2E3YQnWfwgVnXeT2YbtOwVS
AzzF3W42+3NwjqgvOueI9JeyJqIlGLjjniDlkvPdM5iwhJQmT0HFoHjO0+y11fihyxynbW9dvV2I
PwsXRgeBWQizIiAqv8hcA3RjDk1mglNz/vDS3GzRTk/VjytNY3u4JaFqB1RWiJbbO3eHROBE4Nor
Wx5QoHyuLlC3qNNvM5Tk6+CYBBY3J5iRNByOzDH14RF8FYOmUBhJOd1NCSrynm/4c4LiPXhJWi6M
umekRdDu9+xdQ89Eb9eBQo+aPma2LTppT0ZUTDmu6d53U33tl3glEhdReIxnnC3P4N7BItoaPnU/
Il6djEU3j1TQzOVltq4m/1sUsRc9pb5dEFm8Q/sZWZloopOGS4lEv/2DhSiAnwqzAvNfDAPErNY9
MFtj2rVbicasR+8YiOuw1BmaURZAjiSI13fEVarflOlZRPP96H5ahmYIPicNykw8FkfdSM0zMQiH
9vbnN41XM3eTXPBeW5EwG5GzJllSmnZAFOSqKq+A/tj8b8qEBa0fbUgP86Vx43FoBxHp5AX08Bfq
MOPBF1/nsp9ZwjltTyXo0uqCV1OpZzN0Oi2XIRZblOf78EFmhYPZpdiEdS9OUkdlyWXYkS9JdnT8
TI+0aEV4MZuid2/pwoZapW8mKjTJrARz6CQ8fOhv1uL3FZKOftJCxQiFYeJe13hBjCO4tQeNBVTu
gUBLHMjryJwMsSvGeJ7GmPx1IlqTHu8Zt4ElKHaNCyv+a2EZ1+HBVo1/dKTG0opJoGyLDcHC+2dH
WAtxpQsH7bo7eJgMlcFhrxHHvo0QsVhPdN0XTNpDXtO3PRVImZ2q2BvftoF8iFWWBsVYpvLL7mQu
zf73f8rYMEvhw38tC5zQHVybeetna2ETEzpGs5qyJ350PJo5KL0f4XwJNlG1uTGMo3JA47WqxaWR
Ob+cWahGaOz2lcs48nAhqb5599tbLfuvSI8q5rA+uh2PR+14rlEKJuzzuGSjN3+O0gZBgKQxbKsG
dl7zZNR5FF1DB+ilDlU36y7/vtd6QxFx0/4ZjV45MivHYV4qmYRoSI57pOqnG73fIColpdYH/rjv
soFkSVTMy57MfNrDYeWp5jswna5DUjRwrfBqWKUlLWQBK/7bE/72m6fx651lySUw1P5KyV3rnN64
P1iE2rZib1dhE23mSbM4FcBWLvdwIhl/PcjCw9Vl49oy4it/CGau9x7ZFCT4jlpDr+lwUmhCx1cj
2+OaHD4eJ2ODXptT0n8bhnomtd3n6wC68hhA+nUQJSAEQvfCyIOLcv4M2DLHWnQyEK5BsWfJ1JTr
Eh4XP1wmnLSyu4Kyb6gKGnnfXRixQ3fZ3l+VfvZS2lSGdPx3BrQ1pBKJ6u7qITLFW8F92V+XzwOE
o02pFumMcMejQoq5obLq77NJIWmeysykgqwSEjuMbM2GZmf6Ve8+htM97gcXpg4jkej6R1E8rexZ
shxYVhWiiznX7KN22lxzvpFmUordaTvtJWAJwI7B665MZnL4pTxgi8QnFWZuYUvX7JJ92JNId4RT
x1VfSDgvqKZp89HshqTTY8XDkhSVRnq65MB0ruJMETx9U3lGEphnitLV6iEyRmfjEjPOwI2zZcrd
B9YuUh7rfr4qr2q98uEj0vkENLuxLnbaRsMEgtqwne2C/F8Z51VfRXMtoyLWwK3JOPtRGTB/+wRM
Sfl9dAnN6qoXiLxp6aC0Z4mEmQSIAEHAf9oF4x0NoW2mWchXQ2nb3xg7lLFNMpjhjZunzsp/0g9k
Y5cXMXKnRqQH14+lulw7rOliQplOP0wztlY4Tif0br+JRRHLrM65YeCf1lZacTpWmpBIp8cOVT3v
P7DGpASby4fesFRmONy8XMVcZR51+6/7XTemCUMNeV4KuHYlrEwS3Ib5B/FKGq3Sg9BRizESxijY
maHaeLx+RtaFNajwr2/nVeXoUoKLwooz0WhX8rzqjSfLOs6xZ29n1BDEnVg3RoLYAxcPHw8QKg/w
MjpxBvOg7zK0bcwLRxTd2hT/NwSkELx5pnarKUT/mLK9hSkj2lbfbFK1WkyXgwD9Wpnf49ut0lm2
4WSGUWpD1o//XY6dIFdXoi5WNCufpXTAKBeFeUoys6ZJbtEqxxdhlGkblhRjWEmLIgwaAYZjj0wl
6TsMjvgh0qBqIaevsHdO7WpNthpRnw8FIKPuIfLTSIrzhx8T51a7o33C948fSE+GEY9nEFbXpHE7
NpcJ6XUcVyNsWJ6SQTLkYO3LccSvGIAFwic7GN95dLapbRinBbJicYm/ZVK8c/oQndpJ06jDrEPq
1qqQu8WykPWwGiPg9lz8UGKgreNaZkf883APjLhoYNt3rDP7ruvCCa8c7unxaHPkNPAphPhpDGJC
BjhBmx3pwG+2mx8Xb0k+245q+QIkD/rhPlVuLM0nXuD+UBxWYSxXJkAAP6ua17QRlaM3V1J7+Zya
juD1i9ws79U2sNYcZwiaOieC57VKtKaajGZawF0Iw56s7jxKyh1u9T61iV3+2gIgK8hXaX0/c3hA
dgTf//mxsHGIeqRz9QjrJyFFABE/uCFqcDw7KhooVQwE0ceRpWKJrr3RMdipxRAIKJ0KmU/oGvOg
j86fZU9KnjtKWgUhdhpraRIimDYSNv3p2jsuzkq5a75t8OoPf1mJkLPK52x5Wdfavhp0bW29ORTx
a/lBh9P/hnnB05w79BaC1qsa0fOg2ZrUVs5ESs7JesL11s6JuDeqF40KUZbrgjU+fLrcjL4KwIah
+RjaufXqntHN+Snu+I4Si03SIundDF4/lqvykWciEwqYMa1cjE3YDh8BSWcR6bsHXV3rtnlI9ygQ
30tGEl/D6kgyglwy1QHcGZQ5ZufY7IvocZgAKzbOK70mVcMybXnLAd9pLisNoR+xxdBrbKCg5roJ
pptvtL1ds9vSVn1j9ICw8b3FZ8lnuUS8BIf0A5bV3dVrrJ2msY8T0YFNqOjNnOJ57pcIlntCetfU
efDg+X+o27c1jFM44nG/c3sDVUYk0Xm0Mq55Xgqjwpuixrj1nMOfAz2Im0H2N+neeYO+sJA39h3S
tLanGafAF3SiCzTeWhsSXl4Mbv5l68XIUG/rArhnDTFov36nClisH7pOkRP5+Rx1K7kvIqA6JDER
sHwjypUgddXR5nVFCr9rUGv74SmaC3/2pdNM9XONDxFRshmxz9dIAbAI6PExhiGAxFiWgdKLuNnh
CYppHhk6ENsHhjIz4z0tpZZ3PvN0y0n+dDcIhsslGgRY5qvgEvCFWYtHTBCM8sR3RA55kTCzMJPe
q/0H03IjPThhZ4sw0woZbhtps9vySazRpkURgn7eV5UyT1GXYATqwlA82ku9BHsVqQ/17YZu/x9r
8aJBZB8Zb2boKmARCbSRzHQ+feEmpGCfnc7KRtN1Y81eOisn+GpYj9ixns6fwZF6s/55NesOizQm
TzZqw8QEpO2kSnVwRd9xPMTc+VRQeZ4LfrKw7bd0NC9e3JqRyUdiuaFA+aefkgvgBcg+TD8xLhxv
K6p3ACSjLVxQyfx0Rm4okwlUTDBpS8dJ8nqLsRF8NuHBs0/8KSfAnZ/QagmwGoWQoBinGHJOxXYU
pCorYPiZpmAzniB6CEnt2sy7L5suPLXHTCQev+bnHX2SBO6UwFwq3VDyS43dBSLIf9frwQxEJMPn
av6GlYi1gGCMezb5woGEk8Uuf4Sn+9s6h41T8OB/WoAdREG0Rycm9Y/nz4QxINWYxsRhktowMMiT
lS2jcYJir6BVkHDqFeX2wxQabPRB+UnvYt1PBXOpoSNEOSA5yCMEIolwwyaycpv23mVvkXACaymV
sZyzSvN9zuSVMwvgkv5uVB2tBJomXo2uISlaIrVnlATnh/wsdTYY9DLMdC2bhSXCwQ959rdYbNfZ
MANxdcRnZwjWs1laAe8G1zpmTb2NOh7zeR0DsAbkPTxbWDtUEaGSrjkytm19BQjsMTrQsmcvuECo
BCI0p1tbdbi6RZNTQjRVGM2ZWGSETjhy0d/F4ffOgvm9gha1IELHn8asAW2KqxQhr/52K7vk8P2t
96k4ZkSIFICP2YSfxriHQDUfW5AR6sYDmnfiT+iC1H4CbCiQbtHclhNU8zJA/+y4DJEhqYltWH/g
wQcvq1KBcdnBTc5wnpKgOAArGrd2vqBNM7v9IextTJQpZ00UULs52/vVkC6TZ4rMbGJ3ExgzmtIo
kkYg+w78t2DP+ZqQCaZUa2YWNefYViTWznrmXHlMS9nIKF5IpJVX0B8dQ53H0uP0zTYe+PtTeayj
bb+4Pqg/B5Fsy8BCq8zfI75EkeAguNAKQFvuN2T7xdg+K8n0wCMyCmZ0NcEeFZQKxrLj2jzLzHbD
VuDZqVdHKMQd5AtACrZHz7S3fVdqEvRZ55ZzgdZL5Rdt+BVxnbtpL0jlar/ck3FcuuIWOgyNlwiH
RGapV7LI5QsKCNy/lut4iNfD8WHwkeZfpvz8W7ZToKY5iYW4FdES4D8SE2ThWwetIZ77Dxr5wf8T
FuP57c40Zw8emKJ4mJRu7HYU7+GKwAd7ESVzJo+bzXKLRnrhqR2duDKezI/bLOQCHgQCqhV/3BVJ
8J+tUQA9JeZUEW3SmhtIkjWjO0VVPJAK6/2zrEIMG//I7O/6rgFlJcVs/eIYjlhGd0Zxam9fmusX
MtJAqyA3+MUW2DA0XKbeQN5ebJ8JopMIyLnpauVoUsDHlH+DdQ4OnqmQml0h+lnBy1P/rX8lX1zd
ROL6a37ucRKl/PpoWbrgegMcFXmennxy97dPxGOFEdx9mOUd6FaNbKQ6UIS2RTLwXtgmshcH0BSg
zxsucLDLiSwwbinbmI5B9SESSctayfK647PZQXRqvpcE5NzEKZzfmt3cnZqhP5k9kUklYQ+A7uNO
k4uB4v9ws27aDOVoA7MTOVnKmWZ39nmt6zkUh6UHxN6JMQftOo7XwVYd97lbJ3AslX2I5Qh/jjBB
h75NFDtRQ6ZK7xe+vlpSfyBiXWXR3aErHA5Vx2/0QbZa/z7Z6KvXOXyz6bgkISheA479MxbkXvIB
d/PI5Vxe6V6XPtEHOzciXsLMCojfi+WRT235Or/nzz99ALOGIzfEkIrVG/51d7//I0luT5nPt20o
PqYYP5YkflcfPd2pGdODOJuv0NKS9XFOFBH9+RCGnp+s763oZnyfDhRX3zH8WBv/Dxqmkf7SUieq
eXFAu5lA8fWQuLveGsmSq6YUXOQQCNnyxDWO5x6d2FTaEkhUH4dnpxWym9ND5PA203rcyY9PhwiJ
FSGvvILNFN9H+5zw7EZpVZZpBw2la7mWlFskmfyguEYsVlnIY3KXGIKiAfeimMANxU6YkRVJQu60
IkfLP3wstfsHJDBc6ltXB2XnPWuv8LDAQ3ivSIQsdcx2IHYyti7WYg19GnxrcUZDhlWWPZadFYfZ
rk6/8FcnZPQR/u0Ojs2bykUcvME0ufIf0rk6DVITOrobTeGm1J1rGSMGTkEv4Qub3PZ1t97QkZxx
1QR4EMS73xPwMxDAjZunuyjr/fMMH9Ur2GWfn1X72DgZlp6NbrHvd+LQyjQMBVYAjQkFCurRqtUm
99RmB2ZFyz1hbjU9AdxYQn049OQMcyCPrfpEwGUAPyJRcIqIh8/9t9cQpFClGPfixQu9YoW05h0F
aSO8F6Zv1YwZA1Lz7ESWOReN/GlmfCNJXSIZy5UP4/Ctzbmui2qTpKJMryZRan18/aBDAjUxGLeb
n0COHP1NVtEaJnGHjTA4FrcocF71zoQeo+uMGAVKnv0dlprVdJElsKmonjvNI60qofgCn8Gv31G8
hKOELEIak3QnFFGRIur2+A3HojMj9W/VJuiOQGZFJMHzNifH9YvTaVb0sgW4+cqy66AJ4TMT+OzB
TI/kQW2hCWBXeHFF+rzumMF/OdUtDeJHfCoxy1m1cxRkLf0u3pZcnRALpRZ5RKofTtsTXZKwqK3i
j3TMisiYwJ0W11zJa2+x9d8QNZwXGqC8lWECQz/MJ7wUChMw4ZLDe54tHEx92oYR78wjjMqyZ+t4
IDYau9SxPLoUsHW8EjIfG7BGhTd5WYN49qTknWdGfu2+OKkcRzr/iHBJZPVdB6yQJXIulyhVlUwD
Ah1ABn1xrG6ASO1YcEGrmCYOx2vJNSrNy1URf1uWh82IOw4r0WUuGNcaJ7uWaoK4rpc2u+CjivvL
S9AwGAAGeK0bOwCXfZnHoMep9P4qp3OyEBHXnKwhhpxdOOdLjz71PhFsEXgRwSvjKB7H901n5V+d
qfBXbkAmeWh9R9D/k7aJlDh5m6GKkvz/rPp4E+FQ00RlDcpVzUHFGPhuE6oOWIii+XPQIRN8nWOH
VLENW6xLQIO7uN5e/0WRROoYmWxZbcXK1GFYp1GDwx9KHSfUeVt8GUqyx5KaWdIoMkoNfwOPGeJx
T5KffCaHdP3nO52oZYmeP6uuOwxHHdKTlmsSLF8r2sMdOIqiP+1tlWR+QFCOWjpwJQ5/vaF0i28U
5u4/8t4div67GFsclTH6N6cDiQ0+6OIXqMG5Q8z917Ss9y2oCOb/T64ckHv6XvEDX9tmHNVR0seV
nyUOwRPq15cLQMoiXsDQT27HfA+6XvKgVRsrhZ1mclOyGhApTMjeA2oujKXUuXLf2CkXuY3wOJez
nCFhccu25ERH9AUHYgK3way663/4XoNM28vPBnrLvNvA/XAnSaWK2FuJXn3kNs+9mgRqt/d9xfho
7lF1OrEwIUrF9aapfbFs0hCjybNF14rPTWsUa/SvmMGin9xPbWsnWUGv2NJESTmjSJG8KMmsbGKk
LO0rm15v72cN3H21jqvrPYTu4ZYcKf+lFmLc/enst87YbV4IuHnnyrrbYqPHd0mMCY/w2jZsxNOF
zZNYnoSiZBCq0Z5+Q0yhg97w2jjhQk5/7qb8XYWRFzlUix6ICUVhlZDlfScLjzNMY75worPTBTpu
oexAgzqtMSpnUUxZE/a/j+SFNCf8Wr9t07XTxXc7MRksqWhjNmNq6OKOmd5te4ojogEMfFu55o/A
3AgB626NGKg7YrmemjNGPeYQ7TmHxX3OH2A+mE5FHdWeK9jvLTXIWJmCDMo12H7gY2IPUHZjYu4a
oivOmvzov1keOHLE8IBX/AOtJPGgToaIA1ZbcPYau+Cq/Q6IdYwUrvnqNMaZ5p+m4baO0uXIa0hI
QfmFNTTRmRWm0RwVGGTnJqrRYVWpeBuRSyyc/sHrV9208QfUl3FJNzrLuI7cphocOACwdhHPHj93
Cr082jU4NRo8GCt27rh0rlvO9vh7j34V+YypQkNgJCw34QSklsneqA/heaecsL6ZLakjnEmLnBTa
geB4ILgmKuDRFmr7cHlQUm4kaRPVKvmLdbSGmNDX2AM2Xi69Z8B+92vNCWYQUA1dfTrcpZ7aEI70
m4hRJEAWVnNwXiFjmxVTDr30zCMkKl7RKN2jmexo44VBltLc19VBT6bttJRm8aAbFFajsXJLlW+q
tEfZxYquvFCVTBfkU20jy/hra2IZFvX32d86tRH+ApXAKQrIfgfU44k0RDwzgDxmve6O9KZVA4km
M7SNCZWkOwVGPyEFKVq0vfEDiOkTCJfPV9UZee6otjFjaXbQqwf0UBaV6uAbLs7mEGtzY9nFHJvT
RUScZqc6nH8WGcGpVZRA2KcKyFxBFe9utDAry5EgIyx52SpSPCKdiJU/0j8gjgBeDMWBofaMd1pH
Lsu0kCHM+mTXieoyjgo+LAJ44HnjPOLfvyX6SmAsOPFBLqb4Km+9U0SByH7cEX3pUezVR9tWoJYK
8lQcAItf/1RVVrhD98Mg2Z/tBzUpQQNXRhv8AeZWAdXuJXP7CNUDzYOv3m7rHXbTpoSE9PPOJieH
qlIi41AEOfaRsNmKYoe1gAS7Big2SYWlg1R55jiRxhQvr9nrvJDb2RJxiXRVgx3HUUyerB09+9gQ
K94PovCpmEYpw96KvinjJCuuDoNToa2Eyp9v/4lNFplrPGjPHfkSFPJtaMKRjjLF4bRlD5Fi89Df
vJnzr0mMPRi+U1AqGNq+GbaWIJIIvhpjv5GnqREJ8Yt6ABCE6RxDrXUFqp+8RMM6duhS7UwEUNrZ
8hqhEgH94Aj5UPw7/+LFXhf4fGMY7Olb3EKmwA2Gasyrw0rKA2nsk7BMxi21UbQEQZ7j+PbacJAg
1X2bFkVUU2CMVwJ/d9f4sFAOhFhdpMlrswsbBwLGwV9ydQTfa9rllVRBEw87dWkxTVULkgOWKdYz
7hbH/yMn94n7F0Zmzizo6nuF9RG1bSwJ+i/YfA332O6xYWEsadV1nuomKr+eC46oUsVbN8nY5+Pg
raOYVBmKbvkuzXq9ATLCImEwYesUsI0volglKNcjfgjqcW2jsp2bkaMf1RvKQAE441Ni140RBY5c
CLAPjslgxPgnTOf0cjld9rIA3q07vB5UkZW8L+i+NViXL7mBnEr19pGvVpugzv5X0mLSNpFbYOdH
AM7m2DJP0yjsG2cSU0AMgSecMAyGobOjbelz7SdVbcZDUp2MMSIaIqyzI79AQRemCTlwcx720Efa
sfENvzaLSUIwQ0f3gnvRzG9XrwzPg1BCCIsjV6ru3CnztJMKYB2FLOXnc25hDm5rFfLVZ/2Hq8fI
e79QbU8Cf/B0mYl5bvAhnXoueR9cdiPgH7Kn0ylTcdA+XcB4b3jZ4yypb1MRAIOwRAPCmTKpISMW
m1QX5PjD+0ogKTeXE+FeSLox/WtYJYgLJICz0ncqbrVgaB4nvM08/SeIq8bfgN/nB14hK+RC8xi7
8B63ps0+tBCN3IkyvjAuGtl06zdjq7gTvierG+gdfZqktUrF6ZN/AtHURoTZ7bMzo0LR0n/qJNHJ
FAcVVMvT44CiXCKNXCdxC7M9H4/195vdKsoePwET7xocaTbCCS9+FEiTAg8X+pa1o2rzb/XUwuhF
disAfWIRpyGR/itlUUuL88eBDCpx5gVN+Yue0m9fglWAJ17eRMNggxTLBUfdxoJ7f1QEUF7r0wmZ
GzbpJ1D7/mDOQlOvVQheuoy1FArh5Hc/8k74S1ZUYDro75162JCpOhX262CtsMnr+Nlm+6QMiEjw
cm0q+bKI2bwJU2fJAenNDYKr3DT0Hi5F+rlYIX4ANmttciXC8z8NCILaEDSfiy4B0DUvVnyvjqqx
0yLgby+SUDhLJ2CfWFsFQcxXeFhgeHDxK2lnyCLFOZ6/ODXPBvHGdwHj33faZC3+IJPetz46pqUJ
azN2VhYSer3Ly5N57kifQzHvUBXVnSxjBPkJpkzrDjkPpblUv/bGBF8SIxlfavLFMNoi7QNL750Y
epkhiFcDlfP/TJKEBmOJmFmctaaRNnyCWDkXIvx2DryXJmxF7Icu3V97/IHu7R4T9p8t3ySoYaIc
CWho3Wa+6ikII30v2hGqoPJd30AAc068Qb2wqW92b2Q7SJ6MplOBdibWoXBkr5eQ+3zNjgKdciLI
4mj90xYcHMP5gZxCiv7ZxqhHYjQCqqxVaiJKr0B1XYL9TH2PZl7q8OGUi5XlJtykgymtkqTyrLm7
l7+ks0tmarL5b8yNtuCrCOSTKlS4hqu10EC4wIDXRgMSjV6o1Q0fRyPH2s2l+8uYplaypcODDITo
IpPPWI7ATS2/oLBt8iGL3gwdUw2Fplm+XlLRjOev7a4rsMnrer5vDKlLzmmaY/PzetJ0WfERwkAP
DVCU7t3LIWGBLZS2vKqmsmYEWCKp9/ElX7QTEC7Zip3S8YueM0V1A04sGNWk/m7xqJ0ZYKUOz6gA
hAqzROda/J2nUbrrPFsTpUOA7Kx0jqAvm6UezWU1HeAgC+Q8FsyJ/ii75MtiG75YKY/XMoan8NPE
U0ry31pWJ6+Ipjg9oD1dfMIj4QVzcx3vQSo7qoV7IGhWyVh65INWjzxdDlVyxrdn/KOsS4wZjlPE
N4Fs9M46WL3cpK8H/kbIlMINg40jaqygOd4z73ggy7gEp9LN9qp2zCzPXzPUlEkDWN/eR/vCUxaN
gtXsjQto/CpKlE6OLp9Fx26lL29ZFTrmY+cBMgImDIhaQ98IqJDEddr2LRyiomQgW/C0j2YdQcaC
qwnIWgadpf7rhxXk0VIOY141iRL452mjWpU5typkJ1mtXlaab1DdGjig9JX9fno9O6vPBy3gpK8D
YVlePQorAs2uAjhZYXwrLBs6RWBW+hXOfIw/N0IJSQCaoDko9BzbJ5RY6xiUvs/Kk7RKSNs01Eyq
7BQfFlAFuFY0rBO8cDrRPNXinDXcVr7Ja/f4Hv9BlRrA6nJ0whKuopE2XPZ10K4xwFsUZw4Gtkkg
M7Z9cBsvvMgg+gC/RnlbbrcCL7vSK/2x6c1ZtiTjVJuHj+sAprbmzFDc5dpCvDInE71J7ORo3SnN
BBdjY5gIy9ACJ51WQz6MOJG/f9Z89VIyOAx2fi7ZTfkNuRz2b3yEsVAUVgLCh+wAjPj3/oBT2OZy
oHYQekQE/6A429SN8qA+5i/DtoomvJwT4k8l+XyXpOiDKUqyTriZOOkIasn9+0vciZkdC7a+s7Tv
sXxxKAKfIbMcPjiQ6fILEKwTba9wMjbsGoYGIsiMP+dX6kFNNse7q08dYsmBBQRohZZJ9Da2RBds
CM90vAhYpOsjRw2XNN/lF1wMXC6L3v5+hB8ReXtR6xYUq77sfgMAM+qZMUjqHyFwYBW4UY+hn2f6
HRyYw12eZbEH2vxIYqca+v3auCo/kmhdr2bcbHeAGm7T/7E3zQPFjTLXdSFPUY90ZwLJFffc2Ebd
a8D+qkEeqTozMUPJCMlJCBcMUk4wXwXPf1RbLtwYSmumRNob2n4KxKvwNIzgPZrSD5dYgI+thPMa
g3LgtRilSWkXNWOMLc3udrNuU2CtT/CaHMLgNgL+tM29XCIPVnK3OpZ6aVoS5mlAvCBXF6qheBDI
sx8EM/ZmJ6AW3ypc/HoIOjvlajtaQfBKx+j9aSymOEPpqF4CD6GIq4hU93RdjdVgCcQqr+bfLhOO
aELu7nI1ME8mI7IPTdSdiEzG8rhFPn39nr7LF074ujkUAoPv3vJ/xZ7awrSQyk+911kNvst5PcPE
iRAJmC/qTCdDnkIVBkBb1O0A08aBfQ14egkEOgQQAEY464gtWZadpmy5afisuh3xocxIR17F8BUO
wlxaQJ/62b3zDnO8oOkhkpwqWGFLI5QyzRn1iPeFXK+k4G1zpcZWhvpue5HE7aXKTlZuemy+ukJp
fGnitHh4bKEz/RbTdm25DEcn8i5mCU1xsXRxZ2qmEPqxSeiPe5jrsdzmcG8MwJZzSbwM5knqBedl
c33TI8H8aQ4c+lEcM4YLyx3ZnbgSx+KnIE8cb1RSKjwm4DcoWuwrwL8nr5Ov+wTzeVl2ApTyHEe7
LvfR/KmsikGHWpbEaEJyUbBZGUQLja0MuTBXoontEW07BHfRfMxxVOs2AmVfcvvI2FZ2MIK29gEx
9tDAmC36DNi5OLypUBC2Nnp4xSRxE6notA0iVtG7M4AYHSNR4y/BBKst+T3rLXK87QRyEytyfG4v
BxTDc3vZ9nGXgIDkNjFPA808FyIa+UCLkQvnKZYZe72EhJtEQLHJyJnJWkVdjF/u0WbB9zBhDTvT
zybzT5VRGMZxJ/4Pa8jEjGJ5G6us7COWOtepzwDQbiNm651lgOyVVgeDHeZ7IgZnsJVKP2IK25Tn
gX8U63hoxZEOYLYaudrYm2j35xNRwCOX+ig2neQGwwWQfKiw1sj3GIZc//wRad/fqtAOsvsdj8wO
udKwtW9+n8aYle4k2o0XRke52wn7FgllG94J/fiwNNibhMGAtNPNLM9iwD/L0BNicx5SQ0WZvB8o
DS7Qj2o6fD+Oelp+eeYdK4yt24pDgvDBOE5Hyz+7LO9vkYbg6/MzpfQzYhTbSWWAHiJxTcUI68UI
YCVNN8JGgue6CiqlwduCXLJwEljBOXuH6G4lnYEj0eW3WUJvyOl2d1K2DowwxNR1YaLDUn+55acW
T0ggNDtmCheQXYKAqhPuqEIrxag/W+XrOTCbN1t7dL/oHvlYg+Z8x02iwFfyIqNfuGFq4sHLDMzU
E8ABVNWyv+ceJS/OHBhq3S/x3VNnQJlITNWFqef/jK7Nj9riBfdAqqHZnkvgNo1Z9+/TP1qeb33o
C60pIGskKmJ+hkfJ2oiOY5FwKzHMREHfunUp9WSzgo97teFmhWTQdn57ukbbpkVaAWRvK3P80F9+
Lfu9dAqcQvq5zpeUTBz3P9JRj90UKxZeSowgRdqqY4I8xiO5zrXmx6t5Egl6SkV2ZXyJluf5GQEs
Tu7EUOep26WlIpWjwkvz6XDijtUC/2v7zw1cvqJhWk9zMpKahJQrAidLtc/HBnGOiI5iodb2w+kF
rkYZAMJa9pS6OqVSE7WyXQlNuHpcSpyO6CZtCdgTm+6qSNa+REvlptbnt/9U3R/yHeLWYhDs/tEl
b1/gMdOkShyipIbiK57CLgw3+fZzDyWCdNcK8ij7rxF632k+W2Y6FfCpSIKHAh1axLjUmROtav+T
R16aKz4zjcJ0ekXBWQ/TfPvtD0zzqDHRdYkFT/ixWNIiu4gUvrX3uO41uo91GWoDOqZlDVslfGR7
q8KqMaJkSiyaf0zeXLbNIPPmZv1mKlosPvnLsOshPkWdfnF2HEa+mqfuBYUIUsT+YrhIJmjAHCKo
Asx98QfVsWivHXvdsDwMRcTUBXXLNVN0vFhNF7NwtTuZgMvvqEGMJXXfwWrM1coZojvo7BjdmMUW
UQcAPh6aRnUZ4nV9jREZ2WktDheIWDUKOKfL/eygSKawLSo1Qp64bJVPheKLYUWJJZSBTb4uGLYw
XdrdV+8dI2nCY51TC+oXPoW5gx1t816g6TeTKNwiu6Qk9pprYiNZihXdnkb9Hgkozt0hMETKSvfW
Zw3UXJHs2ChSG3U6L6UqOJooP18vigB1hDWq8I3c/WcbrF0PE3cJmOJUUbCM00sdUMn0xhHI3511
jL9sd665531JGV1iwnF5po+Q6d71gG4qNlTtV8r+lUpAfg+BbqQnJvnFBMnojU4nkc4kPQlQ9waT
EH9zG5ImWSPFjhSxlGHR/471DGIKMS5Dc++aN501EmWbR0bh0YPG9jbeo/S2sYvfbEkwzd5r4XIH
z3YrjfSdRWPFdAK7dHSJxeGCGPJGJWUBfOk5+8RFLtbGj3g7xk2SyNTV70aGmUd1OA0RnYG4zy9f
8/ywQ2FMwKqPuZakjwsfVyj3PHXNcR+u6UAuQFfslQJPBQdoNFYbl7bos9eCh6uFzPBh5Aj0s+BX
KFROZwvkAhyoCDukB6jCGfBb0JtnMbSJP4Qw9nuxspl7O22DoADXxI9UE3LLWl0yS1Tsl17L8qNi
KJ1cMYfQ614meAvzMTrOHbqTKpWK+ftlgScshgEKwPTMP3jZ0c+azDAM6pQvELVsRIAtK7zc1zcJ
JkgeMSetnIGrgPAyHwt5KrHbKPsFMiR08rE8MS5aA415gcb/WRGK6JANiEHApvlC05gqLlcQeB+h
mVr2JhP/Zpz3iCPs+ugfporV6SERT1Jpkvb5IzJFedNPkn/RZmxk3ajsURacsADWcf2CD/fRfvws
D7x5h8w1RxHK487a59k8qh0Oz368BCHAT8y7ILJM6FJpjdD7CK3LqOBlurn+68Wyj0apUQ2xZoOH
Fh+re/X7ywthGyDP5fPpJ1AcRqroayXntwrM1/rDGQfP8Cm8Oa5Fmgj0Syozp596dzZFFu1lZpx5
l8lJxpz8p/QPj+DcFCi5vbFMvU+SpPG7JHHFv4uMe+CfIZLXWPMzvMETxvb07FtbJuwoiOF1QbRc
96W6ogDnOmbAHzF+35nKlGq4lOtNhnGdngNHX9nEB7uwtEs9t0WHjHJ2ao3bxQLXQUwcOrgzpK9l
vd120z8/tVLzO87J9xYxLSUW+gORJA6cF6gDqF3V/aiYSOzKT0sKImiJbDhvc2TG6vObXPWMid8m
lX2AXMoaSDyuPDXRcGvhy5QFIiLMozWWtxumZDEoEmTTOXwFhvWuycCprNUCLUYcZvE+LQS94Crk
FC5kx1SdMIxj2ByMjTA4H+jXFiY7V3iDXO54XlqHL29+owL30l4CdKoftt1RP9su9I14wVEhXJvV
VPWcN2CmN1TJa1Iu+NGbN4NOmzTX6k0trJtCQDwzO/VY5ObrTQIW7/Nqii5q7tbBaTHoRRX4O28W
lBf7aQD9zG00qpDXphidVqvx/h7yCPB388GktdMCE0Y4gVfGbkxPKmG+PlcTZW06OMFTVXKtuYlK
T5AiPsEVSCJN8R+SfxwsE3S99Hh1kxA4K42gpuy9wAi6uH25dVGV4UBBj8ldxRXCGzodthKfdSfp
6ZhLCZpXOm+ZRyv8+emVPyGvSu7brD/A9yoj72uqkKHqwW3WJ3BVmp8dlrEcYklCm63aX1tTS+cQ
nAnROUp99iIwMYvItwVsly2WBxtXkIt/WGNPfmnAHtBeg9RfRBuwAt9tKg79EnLZjx/nYXOiHVqd
4QwYCsd2xMuYgd7QG74XfQGSk+YnSHOzFmDsxZ3TeJoCxycBdQ3vyFbE5VsujX64t7NLJNcMVqDc
C5FblBIa/6rhYewtq28wUVDkgrihArJFmXu4JtCTSmt3ROLIyIKrD8pdSPjP2k5yAARkU8nQ9glQ
FSDAYehkNKNYOmmA1pFHtqBtEpOptpxDobz5WbfpgINMuLUSNI8RZMzxTZ6m9fTSwVgxDQHAEIh4
zC5KIXCgczImf8kHwxLDbzZl5mg9Y8ZxdQmaGgrRDMopmURLj7GDidVBAzGRBYg3EicHVf/D/Q8i
gtF6ElYKDURzYXJupPmFRhj7xTTRnfIwu09rX8qZRafH0eUf5aQju6MpH6LWGU8Bs7kH5QVRG9sT
EXOftK07T+IYETG1zcyH1a8JBDQJXDWhXaxV1kI1Jrli/5AamKVhsC6qlAEp7IROYsqLFeEF06Fi
MmxxzDfUDmfRCAziLi9npNq8SssJtWANaPzll/dirVxKTsUp5cNEEkmEcf/0ehQi/CERAI+zcLUw
TcIbQzBwUQDU2f6wKXM5B7/z7/dgJ+34gpoujgAoMUYCVKsXlxNT9cmGacJCrPYIbMmDfuYhvhdx
WOrfxK3xprjl4b3yLewp4LJh8qRpKwtgL6tyWlLE9/dAH1mXENSjAshHbZO973+bhdZiAerw/yvy
oAYn8369tm5HBrfshuOiL/I4Jr2XdVfWUCKtKzd8YYVkgx2tfdCB9flwC8MzB9l7d/jlZC9N3bKn
bUbjG0Q6ZrEUOi5wi8ypap0RTv9EDEJpwKXTvoJPaBMYrEI4Py3WOW+svVBfmZS4tWCdw0B7h5KU
bPHvm9Q0gvkZfnGV5yDQTipdUv0jrxyJq9oyhgKhDB0N2Xsa+c1cvYFbmn8YBO/7gw+dSfhdSWOL
DTmDZ44iXAZH6p8snhHQXcq8NC2lT4NF6+/puutn8m+Cuer5++IcruqWMIQ9NTJEJw6q8kTSfWu0
vtXQQjG0wNZcyrLQU+8v1eBB85wMkD1xZfBNive5NzUx97fFHIhdBmDj7t+gl2iYA+LqgU5BUbi7
Wna5O+qSMYtBuu9aZxE1glyr0U8D7JmmesqY1XPiJIGYuCB3+hTL2eTEt32Oz/56l+63ChmW9Pww
ie1PnrqMYdaC7FRvWkNf7x2Vmw8u48mh6AJytpHhPloEcbPUZp8DkFkgLYj1df8UnFev7N6J+hj2
DFLONA9p3mcMYXpMibjkdxmHcFrbP/eA4UvQxCOd9EUDwr/N8i+HVEhviTFBFRSHxTL9NgvoP/F5
uVgnApPeUTp0i762TtsUkiZro9ghNADUL66ljKY7isDWsT0cWyenW4kfx7rronz0qWfNPS2q+PKb
hL+QeE5Qd9eYXOvOrheHmBMSf2yEuxx7vaamSe7quVPKBeGY8km/6bLgRkScpZNTTQgtq6CAUFu7
ykt6zce6a+lHKAIYOhkOuNd6Qb0MozKdnqvq/rz+eRXEM240icQ5lsC0mntFr8SG36LSGUxY0vWb
Bkgs53JDjuCvpYnhLZKVw+e+fxrJY1mHZmkKSEjKwbjK+CutJg0zI0yqegs+M9UKF1MfV9/jW3Ws
KoVX5882cV3Cd8SxMiNHF3zFmb6XeBT6RBxQP7KPvUEyKcxLGsWSuD7TZzxEIukN2k4tZDlxdoqm
LpHnOuhwJlE7g0J0a2C+rC5hVa/iHnrWt+BLdAo/xaZfP8Nh/EfSkrK+0w7PGjLWdVdGO2IKDQ3v
mSWLAYYNui0tkbNRA9w2X9bx07rCtMldc1ruGGXgOzaIAuWD7eBM3ilhyMkDHSU2KCJzgmgEZeZJ
vbNItd4bWEpV/SAVj6vIITx/ho+2Rdie+SAa7Qs01lvkZTni6kR3pNhRpcUPIkdY/anALRGQKCZ1
zXRJsp9Q8RomuqFf/0FnF0R5cV9IyABclku/pG45g8h4w/WzUPAROUWzrQ3893MbzFT1i3dBVFud
BKBlOaCFrU2njx49/kHAxp2TEj23gXh5ifr43xvYWXBVuCjElyov7tDkn/xzzLK1m+5I6WzH/OsC
9D5TnrZOJMakC/6Tr6/D4k5SkySy5Ocj2W3gYTryTD7ibU5kAjOrA20GWmeY+pLYlDkHAF6XqQ5Y
68OrwJjHnDFi6BBnqPZyuxFF6Qvy8I3G1VgcNDKeS26+uS1iA2NSprAzBDfF5QMli1RS23xCeuGG
I/yFSooFTA1w1DcDrllZ699J9H1azi0bznr0EbOcJAeiMJGCjNJB9w2TdpENjdsUEsJ5IaE/2gNx
CvPsxc4Mduk86H2iCazZ6cvdZyRNissIfJW1SfGv1bBQKX61u73csB35SCCLz/id+sTgpKtah5w5
GV8Zw26A7egK3ORFelUZXanuWC7PjElOwrCveHHAOaXVMX/6bYKXCXF2IJJUX26xHSjPMYz2vUXJ
2vY/pJ2EHtZkPa7W6XEJuFb1Dw2iZ8Wno/zGjIDmmguCYnztJ0Zi6T6KxjVKv8LBO8/CRdokzjku
AtJLIGxoB3Wb1nfXGT+ScU+Ubhzlc84+XadZxY+kwm38iQ3yZMdhMCfWvP9Z+7jowosfZholFiBq
BHOyayvEEANmUHitUCmiZt29S7nHdeod5tDdqI7Vudex2nkvVxlv2H5bp/weNvpoeUni+9wv8cP8
LKrJA0Azo933IyXICwuAhwn0VT5Y//poFgAM3FGd1y2DmcRhcKoaKTKo+4KQ7r0Rt0eZ8HUxJiMi
2z96TpkuDNjNYx/fPdo7pAyPI4juLCisMIoo24QDLPiemHHGsKLfvvEIVfETyGYqQvRfTDwnwsyf
a/u2gZIJ0XcluHs+p4lyCgtrU/KhDRCYIrhdPp6b10uRi03tylj7HFKWweyH47XEumUzx6M9G8Cx
oLuOYNUksJIBsbDa/w4kj15veBw4kaG38cKImLyfxF3ULBavJLTu/1ymb5uRH9uHdG2rzTyt0bId
TW871myig4y2MXEu0YfbSnTbUW/pariaXMX4YvbLl5URSRAzks7xK2mxy9aHp7CVuH/QDDoW3p42
EE1Mhwapeds+2r6Q1FLL/LXOd8Xy3PfEkm+qIMYze0DTnX+xU4n7qjSrIYBzmg1LC0nw5uR6YoNb
X7kP+CX/X6kQIYumH/eYJKAWzK38tbrP8SY0SFKylynAaGTq5rqoWT+NiF/QJA6foWlgPB2tk9AU
BUztDf1UK9HepQWqmuTNFY3pUlmzOZceO1sXUvc8BjaFuc+Nx/cdXR466L11QsnNSq/SQ9daSE15
Xwf23vQv+0Yp9cWy9ro54b2RN7HK1Pjj9SQxQXrQhBMGAldcZTOwfm6aAq1mIyQo1UPJtzpvACrh
q7ZLtPB9FOBrYY1RY7sMEpn6w7xQZ94AwE27p186EdD9Xs0fiAEiPb6S0GVkc74Nd/mmUjdHd7NK
m6sUU3Sl033MQ5UKTs03z/dozpmhY2W+04H3LHk2NmwzPbZtEYeXXWQqU2Ucl4vdx+Ez2FUDZ1Y6
V2xDxWfxoQ/mWQNu1NhX6GQSmx1bpyJI0f/Oevm3Pm728o/CFLuyIuAAcW/7zjiOyxm28kbwFHy6
OUE6tzV66VAlh++Vtq802ASydM/+Y1cnrPi06gmO3TQ2nxpEWfHhm+zZ+kxppNYfx8QluqNab5vS
6im2uJTEd3q9Cng06QjLlF98vC6llM223nHyBATSInIkbpVyc2V9jFVNMrUW5TxjPcrUkeaW4HQG
JfRjfb51HmzMTtupLQOUvP7cpU4jZ5QJPPgIT5HLzazzhStpwAms13EMK5fyAQLXWgux0T+f3mHj
3uqjXlM88f1UITcrtetN+3cBdVGJN9AqtOcRS2mQezFBzR8Gp50GTjAc2dt0Tmdm3foZjLCfRwiU
ofELDTqQSnsWeRcHgRosppSG9dSGfFFfu+q7kFqXm0vdctjEET1sS9JHql9lDTCbeSEV5VX6gGTk
6xZZuLWwgFMr7VD2Ocykjaz1J0HfQldsj8bGNnrj9Y8fiT6grQIP/ptIOr6yY7aChTm12jlCsAJe
52ew2AGb0qS7fPBRP0JYt0tHF+Byx6njNbpyU1oWU8hYb9jdvfBTYWne5JbC2Pr40FhC2HQ6DgeG
0mHqQIGhBYNkwgEe2AmzmcMoBdVKm7mjI5r4VjQoNlyQOGAJpoJ2myXs2Re9ZBynadSbeemFnx4k
DZjG38FRJIjZW4/a10piiSlzPOOKi9TE+QaShCwNgLUo/P9wikUkmqicSy1sF/ZtdEX66D6IUXws
Z3bWEfi9zD7KTDPVV7zMn3wIe+W0yB0IqjqR5c+rWEpen/G6tvIgk5xaR+08Vgw8kOnIIfXq55C0
FDXOw1vSQCOedevU8QOX7kzjouvbSSOXetUJ1aZNqAj5MvjBiXIrxfwhpatwslourxREUgDphGq5
RgYO0AxUY4MBCyRr3K9cIr9QVUzRNscllLxDChW4D3RsPipftuxAwqTrL2wGSioOV2WqTe7Sx1Sp
36jZtob4rc6J2YcegY1ao3+VhhG9un/J1UZ8GK+5SjAj1rJRnbYx3y81qJQBenmlJeqTpEPwbpTS
dJ9bcdWHJoZPtAtItoMm8APLY6AEuGM/t50hajZqkgDqOguzzqEgodxFqf0Wty79aRcvwhgs5fFI
PIwWhiWxQqkELBG8shaEfrsFpYC2m3WiJdgNhAGsVWzE6IZl4T/oTb6wjm+INBuiHIidCCIzvn76
50MwKRwDhI3zOqP4I2B/QM0UKqE9AwGtCOKVAPN1ayTek9BlNDz5LVAneSGXgOi+Tm8IcvSlh3lN
DTZsZBCA0YQzuczMpkve40zabPTNWjIoVBKvRbhTswjBffq6nCuU2oVlT/s3XndjQiVZbQlIxN8P
KjSsTsb1S5KMn0M0BZ/Pf1taD0FKOh4Igi3ZK7JsIaqZN2QGqG/7pMIMTObj17Z/kuznwozg9+fo
2wtXamKo8hmv3TO8EfjKtQ0n6QO5vVAS7vDoTbSdjYivVGzMqOh4sSX10gLcAp/YNx9qqdkDUwDG
5sWMFR83cVIUijqetihOv5kOrewCPHw6YqWPULIHADGvfjZ/qPCk2BajU4zEH/gjn9mhl49mAqWk
Tp2dXDyMFP7+vDcHPYKJoPZtNsfdWxRGcnT491WqdXW2viMXOXy3EqICPtqga0Vpf6/Toj5VExgM
zYElamt7eyjNyX4TX790JuDeEVp3eM5HE7lwKhNWxHzDD2+sa8aauJBeBh7DXH1ux9kVzg8BQSVe
qBqXZ8tf+1dAUEQLlkA/wCEbBIXz9LjGBheMslJsfMlw9g67ztktEzERhUw6nA113xGXst17o6Ie
oB0n4PXsZceigSod/tFN1dcxfwaUGXmeT+5WCLrFrDPt/Iz5W1dPvDN7k4po2tpfCHJc24VNU/KW
F/hB7egZUxJO1nwPyWptMBCDMQON3eUNLVL1hDFo15nJtWt7LMIR7tgzoMQmVROeWM09lCO3uoJs
pHmY9/pICoRaoN3U+ahWOyBTT4uvnTn+HAALOGD2aziQxUrUvpQApF9gSwVSvguEPNxVGqTziMLh
DoXLLaMyE485+lG+ZmTj1R14pmU02gOyank0USgu1CCmKvBbGZvdsZ8JK16gtLT+YNwTh6w+jipL
LPmyt/QLevWi4Sn+N+VbFuEc5TPdBFy+zUrF/nF+hU44/U6281HkScd5xKwGLF+gPpkoCX2CI0du
K4VwYbNZntSHKfWWJSyk3eEPPYaPMwuH66CIqBLxmYD8zWvbhpqsLSQ8GqzwYxswg0ZVlQvuxowQ
JVonTwkGfoZLwwgx+26q11DFMa0cbqYqkrkwYirsP9WItLCgC2IKJhxSqk6JddfUlgQQbdGZL++H
nQ+vqdJTQnkRpjw9/5z3HgldmfERsm3CoeJKjO53tlULosD+RJqKvFhd9Jx1iypaiRAPfk20gf8J
jFHazbFswtvDzlv2kG0opi+kki13Lr0iDu4NmIlu3zTQZ1l5nBHNKKTPXeqEVVHnQjgkusdUQgLn
FEU6sq/JJTRVNjwbrnUJZvepzcJVvB9fwgn2sv//WbWulvY74VubABcQP0EPAmkGhYvNzJPYNgcH
4Munz26DO05MYjr0fYL0h19vkYSr8vzMxvy+W+bpvH04f+lP9hXHNU+qjRquQRjjB4D4cqEexNOS
FuJqzrwhnaIkjrJi2sdRyU29ocFEFGCAE2UiMXVSTzfDqyVduxFskCio+9nLwA5/FKrzLhFxR7QY
kpc3WUZnTMJxPsVyz5+/SxnrhQ4/utWjfYfrlMC6W6+07B+znUoKeLn5TM6aLXNuRS9HPyhm0632
QoRZ5PSvUwW8+lUiefdR3BWjxMIpDafjXN5wOKpF9pK4JZP16nb2AZ/KUnrIlcKUla7XhFO8P8Hs
zn0l86H+XJf2pmS/FiaReO9g57yA/cLP3zqj7iN9DP4nKJI8RPXEvgNP+PCLfW0AjY9Dg/MPCh1a
hMMOtNbyKGgV+BMX9dU013qjQXDDdnLp5PGB3UNi2rJqibksP3bXRwF6iHKJ/LxjCzqDV1+G/cVI
yv69xTNA3ljCu0fiZ83Zhx8AudtP8+4StGPtgSRMlaQadHsN/tIoijl23oMaSqKvdnjwe+xMicPS
Kr7cHXXvWDwAQsT6cHoLP6zRYEhRPWZ86hEgpvy/sKrDv3Oa8zER0dMfzsg1dduZBAmCZzQHE+Zk
I0tBRtOt9MsBay1aYANRW/4GVy+6wAtM2UwYhOM2xfnRfBp8giA6AmNVIjJ3M2J7sYh9iS78rhWJ
gK3v16G2xiHu3wl6kcBbbIzesYjswXDw15ZtK8UipSZOCWmwDjFlpFP7/OJ83SWl1yp4LUgaqNVO
YANcWi5NEVAHav3x4akrEXT1sWi+T98gxqW/BxxrwWEmqQeU6YhZXqqdtuc36GtNNMxy21lMTlGB
HTwBOgkEdnJ0XafRCU2aWLENcDBL/M030lxLB1p0EtflZk3PxHx1awuzmgdJwIyQTIvABTIRUyar
/7OwzPGFhMTroI/0fJ3Fpx2AX5yWje8dC12u25TXD4Ew6mYc45JEw9WTudtUn34dMSvcpr8Q6RAn
EKnbOL7k/vmppEbb+NhkDN3RYXlWosjRsBAFFgSI6gUvvnYVCPARtU80E0Rnc4GAZF/BsPZFt7KS
S9ExXZr+z4dWMlKRWHMuM4p1LtAcSy4Hd/PqHs4M1CzVdUywGBWSftU85dV7J/GWnwLruAvxJxC3
3QrIK9mpO/dpnxrKFz8kki5W8pPgtqWlFiapqzy+bjfN6kE8nwAb2v3AHsJFMehDO8jNiP/rtC0+
qKfW0uS+OHnJy8toQBFzoIGebYuEo/UyLhfXFfx/U2/UwB++hN5FHU8PYYnZM4EyPK3WfGCYBUT4
UA6O537qoPq2ObeTds+GfjXyB/j8V+ZBVNHBthMJy9Ly5JU/d459raE7RfZEnHVgfxr7uDNU4Lrt
xmfYSyDCs1dNMbdHkhSe1v218tqsUaVkc1N7ee3byfXHMO9cJ5yFn9i8iCpDDSLXg2FcYjETKMVa
3AfiNZrg3OZiqao9ra5BxxkOPdBWydJLtnnbXLGGujhumcgh5rWlAKQj1H0FhX9470GXxNy3qaIa
hXCRn9Z59bHH8FLwq5B9ToShgqGAUCPuFCT05/CG4pBPv8SB3zbdqkrNon1msG7LYE168Lurb8f5
G+VPury9s/NTQ1vzamoh2ZhWi6O8PzI7PMrxKfXOH3+AJVNYrbghL3zMfY9Si3sXg7vGMgT9em07
uzSTtL9QdwOxIaJJ6i6qPfUAv6pHSVYLlAHU7FwwLhA3i9f1X+w72H6dRkNVx7dlmoKZDkWemQTe
NzPuiqTOlmdzrYki9qvz4bukF2PxmhJjuxkFLmC1HUpgO6Q+8s4qE94/PiIgaCSXZ0PQB72CQKSv
EhwuQEZDgCknCDJ2eARGKn/kXGlCWYO/4E4IQmrquVjOM5LoO8mDu7q2rRBxFV8X+SedhYe5iDI+
5T/9mn4CxefocgJlIbwiBZmj1uGG0ovQ8LWFOm8Lvo+d3HX1nRTVb9NNOZZtsrvfVx/ukzemYkeq
gJxqAgVTYWwYKIc+UQ2OzIpNrzY723h1XoqShjCQARpTHE8OTzfiAXueO9UKFTZuqJ+rCVmK42h1
6ZyuKOX54XLUhtFLgavtH3BvjNB9iBprfcq5+LFlReMYTi21moZevWKtDMur5E7MhPQnd4cF/1lK
hUIi6TZ70SjincHDZmE5HIorgaMAypLTF0uL18AwYDz05k/nlrLIrqr+HHZAh0iKPoJn/HTuzkx1
IV8najx1/ry1jAKvZP8nFx5tG1Nj1SuLZbHZGdxJGpinTMMTQjrzJdA4vpTRNsFAmdlDpLI7b+kn
3XEx3ki4MvrcRffV3ZaUaacBmImZyPW5fGMFo2uPVEYS8er7dUXVoQbm1OnI944zwj1QpZUuspYQ
x7nDTQ9q91DhLeGZ0CJDZk0n/+KwI934wQ9FFePZuSCkdaSbJui6RGIvnjDnIRgt2OkZLifn1lDX
nRWvtR6KWYhcmQHc8yiPI9jS/wpFrLJGLBmk9wKtXSJ2pl5J/CzwRCfBYUBtvIUVGg1/MWCXV6x0
AAOs8AYX+fJ33KW7KuZQ/k/PHXJffOHFrL6IA4iC94qRjhbgthjilxIvr8yDLqT56t09Xp8C/p7a
i71fA9NqlKOP3Ps83xRuGJrN5MQxuadapODa2wcrPhEPs/Zj9wTmDu7gsAEMzM3o39TIXlM3qh/A
rLMGU+VOxqSnaoeqiylKDRdfCG+AjVt52pCgKMN/77ZqnQJE0jzk4SxBrM+wyCU30ex13eEzbZo2
RZ0hNnUFHpXqt/u8njhPynChcb9wbDQ2Qzcnoyb+IsajKbvwjb3lownJzu0SPvS5yEmnmpiew3i+
clIQT0lCkZKu76Qfqdj+mafidgrQ6H2nbqWPVpEtVxUTXMwyiC3DW1lHEJapnGvjQtZPbKv38ELC
PVV1xWykARWB++bGSZceiJ0eNRkbW0AotPb6sFE9A3SbkERNK3yObDLQGOYB+BOIAYxeQLr7oKnH
B881/s4rfIXmQamz8cri4HJG8Pt+7pPyT1GwK1ZVF8Fjp/Os5Lu/dfV6K1dQhZ/U1K/AICoJ7Vi7
30HpMskgcxXJpq1u+Ph1r2dkKIc4sZxgb7T9uigb+/CgESBjrcjxUQJVocRjS75D5gRm8TgAQSxj
wbJ2t2V14a/Gz5ORV59AQJ+6laOsVriczK6vwJk1JDETbQe15YU4PSotRWDX6wQj2nh7MtfJtQ4C
4ipdKZ7lrw7tuID9pgVK5671jsy5lLuhC3EVuie+7KNXZ8GgOx9jHXdEDM3W6+BdUgtaYQjJBPSg
v3rTQ+nPMqmVOioNtIk3SSgozYA6iTUaJpV5H0+6Rb1K9xVO9X4djmSjfKQNMg+IH5BNdab1HRhx
rtJEyX1QZW15/+SC/6BLaO66TXvBOhBCXxEEBdeQt2Dn3+gFXB6FYrC9NQdc7u70I54O7dKzm9He
8dS6ysWprj4x7zV6mI7asdLpxRjp7elY505wcbaLPei0gfnEZ+K0z4WLzzAKdoP1CBpjxy8xjcjJ
8Iw2XhlRNV+CKAKAFavA5TkpB6Xv4c8qrPN0Civ+ayC5g2km8a3/mNTcFzVpvwk7Zl1J0bnt/4zr
t6qdkSkOJRRfMVBKhXrOmE1u9gf1kz7VQ6Hpe1Ag3rgReUcStloGFk7eW48v+maAACLxT8WoiixB
1nSmCrZnnTkifjjdw9Oa4Fm1ga0EanobSyZufVppqWqkhp41mypuHk8dJma6MZzL9LBgU5cXi9JD
nFg4mObnPRyVrDWPTI8rY9bViTmimCTyew0oxOD5HE86Qm2B3zWN1+X+Tr7C0mz4inWE1CnP5kGo
bJ5xsoU67rHZk3FewXfyXZikcutKdVNPc+ry1xXxdvaEMYrVzhvYjFt0hA9ylD2y6vZRsh8mibA1
sesavquHFXn6ls14r5y1aorkBwShsdpZH4jWaTYDNN+2ZQuNCLZGxDgmbtS8FNlYjso0elAn9D+a
52Oyot8jmNIXeY0W/M7CfnWzjEg1MN5hctNBQ5yltnJsm2lQQmZZLY/Gu2uL/PAqN1MkaJAEhqOm
p5bU9r6AnwnYP5qtb97+Mr/wTHBqBeh+Z9IddV2Nv7dSmgfCQC20fCcRMkOyYFrF2OMfEQhQ8L+u
rBQU8wNEcft/dt1qmBvvcjp5IyaP3ZDZ7HOxNbuAEoGwT+X6GeUZOwreRyeiUM1oYqOAM7Cj2Ocu
wdZkVgYL+F/5MELzaQVtspGw32wP412lPV55pM7W9VRBIg7Yl2Vr/vbP6EGoBH78ECBRPbKNr8O1
pzTK1KMS5Rg4DCZ+3I9cDBxTi3G8TWVHBJPnf7bpFItxpG5KHmHW+EFC3rFP+ue8T5uBl/dVTckL
NiiSZrbP+kJxHFI1FJJ/+BKZDQOTyCJIYsMkr4vmfypLpm7bM6ZCyUKtWRfRG5fTkAcuXKdf9hR2
0B4UcO1/xxvRrrYwLz83uYXjo9AksR1TSCx8lmM1baf5+ZcH87n4eIKBVT+thEob9ivFfcbtur0T
m0Upe/o7WwRJ2wEJiTBNXlgJVhXcYKqVT6fc+/uvLb9UeZw2MpF1ADYT1614/6mzwr+be+T2cVmo
rC3Tx0tb/2g/rXKdg+dbOxNtVhC22snyeJqVlPzg+JUhyEuPv8+INlyuZDUA40qnOfYsjXDErrsW
y2Ob/DcTAGV+Si37GawzeEfFL8VBcME4C8/7Xvei54WQMG0W0QL/qbkNZlRRZtMmgpJIJ2PfU1v/
pb3FBA91F7XPdScyBUXsMXEe4IaOAm64thytuGmo/oRr2RnqLqjqV23UmOrSF3YnIy2TIe8l5gco
8RbPwEqi9RbcPGW8ndtFk4XKUoj6SwWvHOFyMLDlOrIo4b17Y47kI2EvRmi/RkAdT6Xu/gDHDxPy
59i4y2uPT5jBzu0Hpl5nembJsDDb5cyV1yRE5+4oLldDdQPk7X938GBun9F4BOHcuf1Tq1ySIt0b
2rTj091/PEGwDDVg+s4g2z9lWPdYifxi9UujLeFvk5ykP21B8XG6SbntsWtBjJJ/B3GIURV1BPCz
ifEiTTaR7SK8lGFtfbPGiqTpiGWUOK4dflZBU2pp8mX2M5+ypxCS08TYA2GyTO3N9Z2RRWIJ39hO
op795BCxSKn0ufaOB+Mip5OoToJiZaAjTGcHCRFITJ75X18gwR93eBy2UZ6auDkGam6B+H532r/E
RCCbJzY6hTkEAXoUvDUd70K8FsW9u0ESjlA+Z+yuFBOB+qDSYpfQD+a41868FvKDeGruIic6QtY1
UA9UWkUH6A1S51eIVO6rPaWHInGmGAfNb9v/8WuaXKBd3X+whz7MKTqwk2HHjXKYha6Q9tzn4BFT
kT6VIs3SNcQZSoDwyobqnh0Ynfj8/71UMiA0gbLOKfF6G3/JE45wesKRxzBu+UaLORkKj19t6AV6
Rdt1QnNMDFqFpeGfF2Y3nLXdNMMzCwBJvmx1ih4OP/WltY4OrfWdPZknV/5m+EVAkAjy8dttDCVn
HvSfjunfuo4rib56zvgf3P29nLPgseVaEMMpk7HNG17SOONKS99sNqpX93gtdPlburjzs0PS90mI
qfjcTMz7sYltyyuQ5N3xs2PY9s70q21SXIXfE0AWsem3x7++ABfTSBrofJxH6PK3rSnL+JHFe8Qq
Lt7/MJzoCCCNWQ5TV3n2eVNB396v7y687d56p5WJ+2AeiRLG4xilf6I+8xCeJ3lvKNuBf+NK3Mw9
go26dUeockZo303zFaFg18sMUV4zDmBJaqIpSft+E2Gf0Eeyi4lQKJIjvZ96EdlwLK20ilEVUxa/
prZgQmAuEuRVRYxNrHt0KirX8TZxJ9Y/8jpxmxF8VU3o57TRNYIhcNAvz07m5IsFnoI8zglzWKkH
RaonxWkP+BzbqfdejnUOT24kn3euwnvHYM5hqZ5/fF5pgmTZa3ATF3050ZR2tdpoworYfLfH8wxs
TaWw/7pMyv5ykUcqKmIgnibVAAs73pYTisWAQuINhRoyRVjFewXLFA6uLWzrCmS7SB9++o4bc1aA
mxQqIsG9U6iHH+gATf94mRMqBEg+5d4AkfrwwU0nN2E5YRtgpgqy3e+2fOJyqHpeDHki2tX0PVDf
3suFX6ZLRlLOuNGHqWHrdYTQcfdARR26k3nMS7ZLGb6+dVeb8l2B+NPXsn8s8epRWOsYvCehbAjC
oXkGNlXrr/eGkBAzfe6Htl7OXJQXXn6LktF0gv2dlIK2I65OCl36Za0IRBc3L6mck9Eeb4XKC/Mj
ZCsIWGwNVIWuSvov5cvKCn49YB9IodtMUnRmLc5vv1Wz2thgUGdeRnCticOqqDFHDFzqJIt53zjE
dx0c5EkNqdgsCT0ay9LZ4IJpOFb76igZy8+oeQzsIiR6eWWXd3Ia2kG5zFcQziyscjE8SSCgRAxt
dtbppAWEpvfFrhJzfTFDffIxVcpjvN0O7n1HVKOvZMDk8yjeEyVMUNyMOl/fHfNMiHXNeOljpctk
n390jOpWK9I0IEErvIHnA4Yk9n0WH37jbs9J0KDXkqkspC8gJK4CGkNJzQsxpN7kWGtzsCttu9MB
irm6NfDbRYnuko4Rz2+RiaTOXbmKuBjkJlnfXjkDX7O2WLez7Y01ybmYJ0EhC4AakwJMzoI2/itQ
PHiJ6mgnwa8S5LQE3YVxOImb2jKaFacPAgT3HE6Sy2c3kiERR3nJfq1xz0Yz++1nAuFUiYwAxlii
p0K/5sl6nHIJuRxYYAjGjuBOOP7fFOW2yCwqot/m/u/xYxGoROkCSpUD6n2Q4pnLbhZ9paXWg5le
6vUEFrVx5f/7InJoZKigQr9VXoSQOYcNd9H6mRTLEzmxCMU3kSWNBLF3JlzWxItfShwRtYi/Sv2p
ytvNu5guH6O4QlFjtO3LMai40DsRbgWDeHffsCbdebR8lh0cAQ5ouWZm0lDIpTvGXfHIemOchc4F
G8Bqas4hWe1ESDE5LSMewaaLZdAyIl+jPnXp7OpybvL4xvk9blvOrNZsQ6xnpirS7VG4cJw6j6j/
auWaXibYQFF9m3ThWR2FOOcxQK+vYfIXJqvXTdMxUIXRBW0b6hRj64FQNRpRK7kUJSClmJsiUHeJ
63G7txIrRuDGdpJDeRtrYtlPbfyghqQcPq6+J9ziFBu4LaGKL0V67uihY3T4O45EEFxaJbKuoSIi
fqchgvFsvuzRvpeGXnBEGfSdx+XCQJGStP42pmCSU3S0shuIEJHwNEZdkh8E2EP7wmAuOVDmynpU
Zh4dhsUlgMok0JZpX1Q7JzH5suOd47p8xAvmH/6YDjsQBG2TSdK5Gvp6JxRgDlLRZ+z94aTA7S5t
PXHabuLjosXqr5c39ZKJB4OYk9xawEF9vshCI/3cjM0J28cTkrTLCFHl1TB9uRBHuTA3NfmbgbvW
oe80jSQL9V22y7jSPpas7Eb9jGNXHlbj2owF6w5XJ9XAQthjjw3l1FeSGHdw3SShc8W0/Cxj73+8
iigiw0S4nb5Wc7P/NycIkwjtWLJmW3PCmxMQ3g1Ng0NZhcT3Ym3u9kMaE0iVfv3kLsCbkztbRSs+
+5ZlyEjLgd12MrMFTSTUTPg4L+/hRLH49rSfEGKjwk2B0r2GD+yoxyQjFwnPVyW1M4CJQ42qg3ox
bYeQeiNam/JoL2ZJRayZoKSda0O0UfJlxO58hzll94ysj5mQGfNPNvxlIW7eZhft9AHUc5YbXg85
KCcN8VBMIWozQ5R38GKLTVrQv7EcYOBBFYfn7iD3nGTsVgGR77P+NSMpZi31SOPfQVOTe5zf2Kii
Airx6XWTmh2jhDIbta6BswBbdW/xT9yvD16+P/9eE29/8ylK3CUg6NL6jwERkEPDUKaAQ9I0yu3h
hW7NLIClQ0tCaM39kVdmsGuj73uJ61sXVvx6Md8RBa5iBljVVRDyOjnicE3RuiQKS8NUHY2WsBUW
FVDfWmjV+o+n24CkoG32gRN05Q5bJrii9/mgOK/fuPkyqgsw+notYv92k9IAKjXVQgTFtNUOpajd
2uIHXFkZ1zyCYSoVxjBv3noSO+IECZZfsP0w1B4ZUa/TFUp286ZtDrUpHiYWJWNPsZeDZBOb0Sds
f38bU86gYN9tka5L1ntoK3OLJW6/WZX6/qxqrhcwX1TfwQvVrLgQFKOm9VFGuYc36bbvMbdyQon7
V9z2/vCeRA7TQkC3/LKLOGequB3ca/GA2wLPArurTXXlr0YC1OKOHolraJP4moDCcbzcj40e0WcC
gWHHAhXKa2tMBcBnRaIupjC7ND8HmXYcEm1y4Qkc1sUrt0In0h6kDmyEHTKtGpHrJsVe1mYQDGfA
vhErw2iU+FhiQPAmPvA7wfc8pNqwTZKKlDP8BNZOl0f4O+jScucwAP0lBbTwyZtIVEV2JQIK75MC
I4uom31TTx+rW5IhxK4xt0QXxD4zEJ7la5RxZDHbk+Mdg8OjmOjtfbCx1XIRuBIP3i3WpAcQZ4dE
3y66I2DvwYaRpCZpEF6k9VLFfY9KXsGrLPfoM0Zi7yczrF9bCj4gDYJrN0bLbtvz0tVsHfTlnLqP
U21CkIeVHdFzyD9ak7Le+dV5CuBGmD/wesHbpcT6mv/Dl54oAaPhZ3hZ0G4NejK17VqQIcDNYbUB
gKke8NBRZQiLkpMYDaneUlM3cUKpzAZLKYW5PHLyqOtxehmTVo2tscrkkLXbrcimTwS1PenUHkCF
Tm9cTc2cQckWi+iObaJMUIdBuEp0T4acSp0Y0X/Bu2T0uV5K9cp+pFGGNhecVcwEtHjoWoSTgr/4
/ngs65k3wDbVQLLPgBuuduNf7NekIu96a0zptzMLZ/BdJPf0vzhV7beiHsfWmUTRkEuK4skjZjWH
LHg31hwQRZWTTuHzdpeiVkaZMmUJ5213H9CfSQjW6bc8ShRgzIBPjjAedtrZ93ccOVwPVjjZ3MYB
ILTI4lD+HpOKvL8TEcFOw+0ZAlOUDpQZ6pYXR5YUYLepydLf7LZQ3oQqwJQOGDbXC725DLxYIPjK
qkw0GD1YF1tKiOD5lhrppdiGPyDOYC3Na7kt72ifGdf0mSrVKQocHVItIkKPsEkaVCdBD/swXu3T
UzC5dkQodIbu1vyo2J+CpkscX+j7KFp8uf3i5/QcqNZQ+VWlQ3YWGswtCkoJ1tOM+wdK7iCuGpW1
zYRqNXXduN9OYMx8nkMAfII9QTRKmG7+Vhpe+6Lv2N6MepSLHFLxgKzT4Qn8LFvI66aFdElEOBdJ
qL3+bp1iD/B0SUjt+VVQGUqHN6JOo1UgVX46AHOPGu6FapQrt9Gk3IKGPwUVC53M+Og55cUruLVc
8FbKyTSw1NgdgCona5l05gBfEqmU24OSGZ0KDtZk7zuUr38udtKAd4cWUEr3vIbiSE0uenH62uZC
Eo46/NZUYXTM8Zg622B7vh5cdKRqnphKy+afTolU1w55MpbxzLcE+T1YdnQ7Myqmk7DUM3c9uMXh
67DFsJfEereF3zRWyAvQFWoVvyNDgN0ijLi+z4eVVG+r0upqAWInbHznah17BzWHwi9sNXdixseh
zt+vgyE0CjdcdkFvNSI91C4bz87d+mrRl8BXk6wCBBOPwNTBnqLUs0mlGH3D4BZJD3pdFS/bfSx5
sdjYHUwsQ3Mhcf4gYzw3DED3Re7aq8VYR0d3cMNs6G8DC6LSrvQnrY4Flz22OsOb6rgtQjev8jdF
x729EevmxKoKqYqNaGkQQeKAXeb+TEBv/XTrqsjpxmUOO/IBpaOpYPH+fRoeGpXWvIgrgRdpmDgD
a1lShsfKZpp/qSctCtPwVQSgWEMhomNHDxy7WLchkZ/Dbkuk8jatUNhbYPwm2pJilP5o1VGcETxt
pY2Q11t82n91X482bBfe368Pu+N4zN6DTdWpV0hfaQM4IiFRqLO2vU6XNfkNdAsW+XLAYw9QvT/E
9CaghQ/5APx2O5W+UBejWfuDsUK+uW8Yg60U6izc4sHUP9eX6+PzHf/ghpnjxe3iTwV83KWinskQ
8Ti+KJGl2ljJMN7KQq6Yt5Xyi3+uKfcgG3Amvqtj8D0SqB+r8YUti8ItiK+roWpCH8p7AKSng0jm
jf1bTGcQV4+ibbIEUQhjFeJ6MI8COfjl0uOw2+AdQiUVu4WkDjqb5PLBP5YMfTLfkD5n6VukVxtw
e6WNIYezc/nFuyDzgMpgtvXLOjpBILa0bCsAfj2YlG638qd8kp+v2bAjSHj0oXR2wEhsSEDs5CaP
gLSpuBV5nlJa+ItZbFk0l3YKabA/Qtyap69V/QP2ac3qjP77pl2kdpQ6rnj6BuZlWlETG0M4AnF7
ofNL3Uehn+6Rs1KxxGL/h+5sDj2exRufdZGzni3GQF7LQ067ZG1LAaqqyrhNRGsj3n/O8ko9fcyF
Cjz905OsUgy1BWNja+jSi6DU03K8jzJhVcE7rzU6TaX7O5Gsjqj++VG3W0z6BwGdWODxUAdVEmey
GRJ06cCEDtZqvqaWBac1jVWCMYg98r6FQL0QOYt/nZiMdwaWXiQU89hJgzaV6zL8mjgPdG6uBGEF
7Oisx28My70z7OcIjn/AYdMUiIIcyY79LvZyF/LCzM5sxFP8pafX0zw1fTV3R+CwRU/Sv05i994f
k11YomNIn9Q3bycCSl43p0ffNpXE6LiBu7GEaKpuc0j3W802mljeTyEptDZv7rMOj9QUe4DQkiek
Xx8UbH4fLn/L7+J/nLJVxTNiovHnZxLCp1MwJ4ioET5VtJ3x0Y0DlAuBJ9Zxs1KEXVfc0PT/HzB/
GS6s6YCKvXanPUk/K40kXCllUGLpPR/gE84pN0N68GtTDjM2+2CGUpZFhUwmtGbG+AkM4NUpMgwj
lfLew6xLLl+j1IXDaPSsy/CKT2WKoPfKI/ABJrmIopvOrajX9FomaHrPMoi+ytSZOobjc3oW2YTf
G+GLf5aU3HkIs7wtaK+1r5ED8gbQt7Zmomr5EIzMRfRaX9vpo59ytTjpFkqa6PKgkzjQV6GpTVa3
OssSwUK7rHoT0bcImEHjqnp1N0Rkx9cOfkTzgVHImxrCLv6yynqyhRCB0GenDvEokYbZdSRxfrPC
3SxOK29l1XENHfJV+2Rwz85qy6hCI3pFTIZjUh6uks+qxIND0BSWSqaLvDgkC9m5YFJcr9oxESHi
IRlGz3JIzu4A3Nq+MFTCVFyRZoEHiRSNBjCWezvN8tVnMK0C80IS6Pqd5SaW3qPJmj+p36SWtJoj
WOwVSpPq+bK9hedhjmzLAvRrhdgengJupAjbapysICyhxmLoTc6MmN+rr2SEkCDKu6esSqw3Oeht
tXv7WDFC0hScO0jlLFBpuz6hPaRBC7WaTJd4gtqDZYXdOGYF8l/YY+ek2vKIJtvC40AuXv+t5jCP
bO0vcyrPSGt89IluMvUPrjVgCogb4uVcFjbTv/fqX1EQzsEiqTYlvwOEIPVlDHfDMoa20pPJu8aN
VGtDPhasVG05ZYkAvT7QPIcsPSqOc9gBaY2VEvUMPRv/6DFwtcxd+gVRsWIOZ9eKhd/MCsMw0NyC
hJ6jPVOLe+590UTKsYEQRKflENCQ4+LXJsrztG7nwOzNAX2QX5Fa4zu7SvEqnlJUgfswx9WblQFq
+HivHPDMBLjJBHn4heZ7VoxSutFGHsmNinzS7Hf/vjEeH0va4WbnsSkzL6wZfHH5jj4lLbv43Cx2
QtPTH2giQGq2lhgZWgppDrNsTMm9V8vbedcn2SHfmW/8rWadjya6tggraWCPGtUxR2OLHKYc2VSv
40dgfNBmOtQaNH1z6ssF8twu5Rykf6ZH5wMPU+OBt28c4yuFrPhjt0eS9iavx1Wgmr7pGEGGTWVM
GxUhgKiyKPJjdMDDVCc8VpHSlMqcSc5YPqlXPUfADPAbYFjWA3xPoQzHhL45GSOx5RLyyNgRHVNU
ngSbthGQz+5wMAqfRFzmtbFRh6Y9YO4aDRHHEwlm/r7zCow8Zb7yH76A+Ijwt1Tc7dq5jE7I4yNW
E0gPYVadLGoUtLzT0yKSw/dJQIz8Q3bcqfuscU4kdHBe4a/JfSyXkAiRQ4/X5DSuCsSzqzh6Tj5F
4ud/GAGk/PmHPoSirCIXMA8JLpQmn05bKQogCWKdCBkcjMPNUsTVFmucYYDStDNvgrBXMNIwfJk/
RCxQA1yXaOZS9K9eQq4Irop3oZvgEGSulprZEymRD1u55oVCo0fFKGaKGjEmn7sZzo2wOuFQMVl6
VOCvJHG5Bd4jPfRTTvAfqkPoETSDwyZf/mDHPE9MvciLVQSMkEgAWiMKsmhmjA2++ThkdEMIa/Sl
IND2r9zAwkwHsxcwqRAiKPhciMBkpn/tW60eGhxciI5AW0uY5lowAPLhD3X1izX9XErY3HpLZkG5
C20Ps3aEu/9C3CT2KrLHmKi5QgJUM9TVi2B/6bHFi5gD9gqj+oGe6ymrB+BCQ6BKygP1ELZbaG6n
MU8SVP//gK0z/My99o49XiO3BOh2E5wRdq/NHKTGzc4NowstT2+qcQdS5fLspmDbOuTpVb0x0Km+
D60WkSqfXNKKu8FJt7TcYYnWtsf7dbINp7yJubAvp+HSc33Gt90uX/SXO/EV0G3OWCKtG53CjE1q
eDf2dMsWDsPVFlJ3gKbpQm2yLsnmydmFifQImlmv6RI91tsbpbo7Jb8Mx+Jn3BFm+3NhD/feMWN4
k14WuPgHz6ge+Pq8SlI2c5jOIoV5UsotdAhx2L7z11a7TTfDm7rFzOhcTqRyC+IJei29zJ9kXcPc
2KmZgh6Qg4Hoax2sJVXwvp88cdEtdt3Bc7VbphMi4h1x+wXuG1IRsu6GJDjYYgQuZ8IODkUB/fq3
mPqdHl8C654YcLbqVvnT++PPJUzVkCEhTNg8YF+216uuqlPBKmOPuFi3gY3MKtoTh80sMbK6bTAf
EmnHtVB6DohCBxV/SoyoC81lQlr06lRusKf5CdVqXuhqi9j7gtRkgMT6D/CmlJBSSyQGTuubTOJc
EGonOvyvQfkpA+ZkGdAFJPj4Wy5Yp1N3oRrqRnk0AnX9zv2ju3vfgf7nDXMMludzH4PBb+YQk0NH
LX/2/sNoAYr/aG2k84YXF10vKwwn3LK8K8hy+dqgai8FhH0a9TzPw72qVahMZsG2iz5QWHsHcsw0
gKN/cfyYGVEi7BNWA8KpDW88MoOOidotqRkSJnXtiQE1jMOLzyN7tlj7wnfa5ziL6A631FCxKdtS
k/hN98/XBuVMbt0IUymBBuyRqrPMKIH2slxV1iR+0slx3n2P021SC+B4s7LiEUacmJw9KxFaSzYn
eQKKIh1hINjaTsuD4Fm6u434TSZ3tmKyJVTa3S7X2wfr2s76dlP6qwaj9bZu54Dzd7gniTBofPEn
d8OTWlEA30GwFSdEIh8M49zr38DT7CRmKHQf6PEA+dUqjNDPhPR++U8FBdlWxCJvqQkSBfvUBU8J
nV6oMHLTKQVeRuHpT4pm1mQTaME9cck4Jdk9QqpQUCqmD5GGpVm9wdlVZHFu1kG6lVGqcipjmUIS
c0eLLM+Ohx7S+D7D4iVmnnw0nA1xXEw+OddeYnY/lOoGoz9Rc6smHerinRprOXe+50cK1fkpAP/E
Gr4/ZSjesSUx1RIL4djmjAna3pCpGmihVFgzQ/lT+7aRTpg3V2DvKwAUx38RsJGwJ0cPPmQyrMvm
q00pE1dc48D6iTrcHFDy3znRtRYH88MqDueQFenjI34GK/sbhNSI+jxB+x+HT2nGtEIodFwL0ktY
89x9mQ4MiyDcNKd5TWqgS3m45FTBmUz4kxby2RXoet/6LLFWTetS698bejVSWQtk4cm5RQhzP5Q4
yrP+Hu2VBs93U5LA/wVh3equ6PzYnGrynt6RGEbYoIX76wfn9hfN40pa0maiR7cS5XTf1WOD5xjr
5Ts1Q2rCC4cKDP+e6i3zNfNdgBloaPfvBT1Wqj6P8d5As9ct5dXP3AzDxxBn85gtBf1RjquNf2BS
ZgSHH4x8u2auYtzlR5vkvx28I/j03V+RKGid7/uQ14AlJIU5TWv8vS5097f5GgrAD6wEdNUEQFqW
fNV3QyMqT+apzgjvKYh4edet4vWG/PaGNkieWy4eu2yTceD/VaV3jvrMpzWmYeeSl/5ag99UQMb2
in5oe5V43eRpthomJU11AsN4evRS51id83FbfxJRx26INXe3o1RU23Oklwvr9q9jYCRxw3p42ngi
lU11GXIEtYsgGWMgT8DehA8yMd5yUQ/8PmCRob3qgo5JYguzAjUSJSXRiOOW+KwGH2ZZVJj20YeA
GE43+iJHKUNIXxIawiuZ0Br+LgnYYkQ8tUYP1j2ycOaLIb5bgaNQsqAbvkCeyeY1dbv6ho3ScBqQ
PBgUVsRrUTYcMT/1NpXfmydTVNjP+Cm5oH9OWS5I5Wed4hCWr8j78eKzAUFNiZAx5a8++bKm7yM1
Uh1XOa2I8hKKlMjj0pMRLR73YTrVdzaPYUrz/K1hqy/1lwZDgSCDB0b0vPkshvhSJAqowGgE2JA/
ZkzS3Y0IhlfOz56IsVPX6yB7fQMrSQHkdnI51eEec4ouvP1I8l+GKy18zBJEZM4YlQi4/DdfO7OD
rEUH1eJ8Y566NxvV56IBz1eQzpVApKpeNOUAoUMk+L1BTI1GJ5Y2b6uG/WoeCpi1OqLV19QRJNSl
ME5hGST0h4lJAl5QKDYp0SHUx6g2HgjQm5yUlYoeBy3JY5Uz0xgrc5S2hoL4FXTpFimteK4P0VWI
EokhVVidyEEoQJXUYkTmuHlY/zyitPwI39d8rGY46R74jq+1XwoMzCGRPI/JSbzJ3MwhxF50eGCy
mF3ka3gAq66K6VAdGc4VotmhAU+wXQCkHVeVp40CU576sqywAmnkQtHx/veV111YV0ohtoNfc4QB
M1CdvH90B4XXqSW1vtx+NCllye1o8bGSrnKGlPE/SBFng1d5WMfvsxk3r9FzEA1yaXjpleOq/HRe
fECMI84xkZe3zGs6GBEjmJlJ6v8WzHYvZpnWcLAmUuNwJuYTJZKeZLim3LjH2KgU1F8lEzHiyiOi
fDkX6BSFR61hYKF7/kN8zlWLmuAEzTpc9eAODWzMysX00d6FcCJbdr/Xb2foklVZxQoIHfQs594r
xmukTEdVo7IH34foOjLNfVq2IOKBmrKIhiTT/oHF9O8Go7Me7cwsuzryQ6YD1I3uhtOEoWC9s+pt
JJD7BSvWx4wTIzgfHkkrfqptE3OX8MIrLDVFFddA3Mdi5zDF3xaPeiFzKL56Pit+aqTO4QyZjcEY
3n7feEcVukWKC6hbNb9vDehKi3GR/+ISUgOP8X9Kb8973IRfWu0h4hlR1rbcTrWiZ4wmN6N8fD0/
QTLJ5gDstj+QQG2nmUfQGRMYDv9iHYem8KhQ8P7IYMiazfyEk4jH7xfLg8RdRV6d8vS0ClbLX6Jl
7TidPSp56jLHHHoKHMeGtthFtGORbQcokT3yLXeo5pp6+qzBp5EPh4sVABM9m4t6ohz9iC6XSU/o
OZEEZONuY76GaBiJrTMk9co7OJSBYaGfXAVZdDGFdw48BwDVW00Ao5vm5WkJqJ6oXnmkcgIfzM6s
EwCCSlk5b8FAefXWSeXlwXNoTzKK7m0KuTWLmZXHKXcqHGKIEDO+OiBKDXvPAET+pXAHLryza5IL
PZbMOmLmvNGzJE/+1oyka6Qq+2ZaDUSFvw6b6+1GKS5F8rMo9h6jQg7HCklNhJHLSgaik0exMy54
GW/ORdvPDmZkKYymMY0AFuST3p+n0FsRzJijypO8sNMuysvRU7L6FIw12qUuL2PWkxWbf00ggotl
PJj7QoIkV96PeP3N934FzeRYjFAt626WRPefr90MkWcBEsA7daOlNw3Y2OURjzruaZoFHPnolhym
7SDmQ3KXnJZa2ukjwADBJcf+XN1OG7WflyN8YtW2lj5FfHatwpRzEr8Zoa7iRd6DoyUV2BUWK5a4
iUaX2Utq+wmXTsnWGj8uCmvZ1WujKATyCPneHKgn+BZrPhvDUloL9LRl4EnicZwkjkJjgiH2xjYw
ZJo+pymwZ8UjZhXLUlmzLvzsrP7L74PG6W7R+1c+o/BCHi6ec9fkg9w5bVrVIMkPVXfx+vHo1y5n
z4sYSeQwAXlbzM0pd9b5gJgjgX9C7wCVrqJUrfTc4PwTBh8F5TBwNmf+mnqOR3+Wirts6wPj+kCX
rHYE6hpEl200e+lptnKdwqb53RxPeuBRZA039OCj7mtojjitRX4XULiduLrY0Ck7LsIa8WSOE6Rj
MjebP9UVxNVFcFFOJt648ibfOUWUNM5H6dJsX/pVNNHiApYLGIpyzolh1TEyYLK2h1tgdfHfwM2V
qSGVwfHyn5IEejj37vj3plNYwoHc2i++YhFsfe8W2YhFicPKTeGz4Sl+j6Smr0jgD2UsxKn6fFkx
6xvbveuCqXvQE/TjztNJIYQeP8pzO+PZvAtwmZmS7PltvJ0ZtFQHs5d7zpIrQFw3a8zHdBmEoMvT
Xi2OabhCG4dCGkmMbAzbRGpaG1Qo6kEloTSr9adDAculSgb+GqnuP09av0q7br249Dybp2aMSPpt
sk69zlldU5UhFz+VwPAwoi9Juc4e071Lww3dIFCpjONF7qRPceS7JxQgojjZ05Hm/0bBk0uWRueC
ZXombHj87T5RypZCgY4dP/d8bbep3MMP6zgEKlvfHZSmbVScC/yqG1ZjSbY6lOhWMkeX4gE4X2uO
G1aSFNQTzTdzaymyx1SrOaczAyEuPXn9SzcRlciH6qcKXzRWX5igf1k370OcOp6ZOieAkgKstkbA
KRpfgeHKWcHp6iYsw9DmaLBVpDRjKuy/MkRK45/Nakg1Eauxm0qgDm7C1bRgCtlmNxAZWqMyYAJr
R7xbzexY5i+DmJqgalJDMFGVoaWtemAUkjX7bIO1J9RGE2vv7//dGgjGkEDeIJmujVZ3RtvvLA8b
94L4D4/O1TV0pom/Ut70UKG26J/d0XWvw5La23XZ2i2cLFxm5qAYD7U2mUs/lwHEFPN4jxBsYrBR
bJhb2XutB822P0f3VANTAgA1X7WUfHx8uLzvfFudKT3AkfHPLn7Emz2EKse4kOpEfQFz7S37gp6i
ndlcAoXJc3NNqiTn3kaoL1KFpek6NA7N/URG7Aj9GyyE61pY4pHc7OkrCUkfoJiwmdDEs+vNIJ/k
Qpr15MPr1U15epN2Bd8g74CgSmwv5TL1CO9DseKzwDhAl8OH1bqrB0DV3yQGCZyiOYGGXcVnkqXF
bUMA6S75HwnrILODz9BI1HzWU6gXpaSw94w9X399q8WLxzKCQLoqJ9SK6Jxv9fdjxJdBMCAdKE4o
x4cJ0sTnZpOKX1cnZVNinC0waHMWcE99EmLTWgp+RllAW+FZvZem+MABMJFelGtrHq09BCXihmh0
oZhMIcGhlM994FaZtEqZAop7XlcW+0BKpV5qZ94D63NmeAJWLUiyv5Pre/J104bFU1NLd94BG6Sg
zws5OUIbZ7H4XhPm1ZB44FOnktgbOb+YgKbtMtMSESGdi5YnnQtRHWRo+pEpU6bljvghYaHWohIP
CkDIr41iKGlIzs1qkr0EFf9rD6aALx8PnmUUidLh4GcF7ea47sS4p48TQIbayNTJzicnHHGJXfGu
UHy6FvZXIp67L+beKbcrZDQpSKmzpiPnVmcpI61vnn1zkhRnC/Xx/YWCKxw5F4aMcGG6ZAl7zV7x
GiHqQx2b4/dtEUT6orwAsF2+DxAqA1Gf18GQ+1Apt1FKsdPqMyQCA3aoC2/RLWBVPM4ZzJpN9JYC
ExSHIn5uvtepmuHZ2eKvLfCRWDH5EpAbsJlWranc3qwK930DR4B3HjJ+whGJEBbpXAKVWt8woSxt
y6O1Ifsaf79iy1LbIafTaRcLOkdXcYDeRtgfqvQ9DUMOdu1XFHnlFPGgdlpZTgh5FnjLxusUEYpT
R5Hyz7Kw0h5UtlRsiwcCL3BY627Gh4IbyEAJqpTdys9zFd0H0/w/lbTX8f4V3tL3/CfQGeMakRqR
BrlIOn0xuxjfgdAiiVnmdCOwznsT41uWrbBbv5EWUXq8dkgsGD1zaBTooKQtJZnt6OYJBZnclm8V
2AzqsThVsKO9xymBHObdqG5MYL+0ev9Qkn0KDGaf4QIGL6r1tJsS9mHYHtJNWGo9wJVcFP7pFyrq
2E7u+Yp6owvgHv9QHTgzmgdE49u1os+sJiVWBmXPuUqDU220WCJFV0d9p74kWlIEYWyXpOKqhuGn
Q6q3zx9ZmdbcGnAKjtzNqKM+2fXtT5TKg5SPAwtUQ2ozYjaGe4W2tzBCvIo6tEJjPXO/W35mfoxu
cnCcxRwFCoghTxFCta9JV90qgycK0y8Zl2xFF51BDjHRKuqZhg0eI/fCyOy2eKL5xZvu131S0jFJ
7TlHlYC8rVtbSAs3JNox2CgDqaSkOennUcjdV7ZDGyaHILU08sk0f8B6Bak3Utq6H8mefi408iwn
upKXDSAddvIYdFS5cEs/pt+8L0FcG2rSRxGzkr216f9gZTi+3mEvk5B0vGeFJKWTU3WE2AuYIJOl
cgleHTBPMHvTRsjZM47nqkLCZ12JOk0Nsv3thKaGLhFemsCLOlQuAt9IFmOrlQwLbsrse6nQ6RnN
eHzwypZ98WoETmPQuqaPgNAKLTi0QSAKLMejuna6G58UzeeWk3DUmBYcC62GLYV2pYh2x/XgL0on
QBWpe1UI9NttSolmQCUN7BtXzBz2FR+h1SaSnzPgdWeWr9gxitq+dBmAB8AwYngsghiJ9mzGz5bF
xkxBexBGKcgsLD09XXew1htxQ2xfyB6eDKkfrK4p1j+T0ff82ONC59SX6sa8aYbrEUJLW4FEvS/W
n351FHltg1arZEZq8Vtz1vJTMne/7E3bpfXVP9orai7SuIrj3uGWuZX6iLBOmFGO0uShaFF3/N6h
ZarNGXxdq94F5foGoycRuY8igPrr1v0Hs/BglXw12HZGPfHTgzEwBW+jmJKC1ld6IzgKN49S4Ulf
mniCRCwl6O4wx0PZdwT7k8a9cHPPwBJfEEJQNuFSODH6nPdKSSDHtPCcknh3/q/StfEVfWwbCEs1
NBgp6uWaQb9QMyLEnyCo2GWjzsl3jVrgzzZzx0vCHxFI0pioPtbAxbB7KC661gAbprpirMX6BDhd
ONeKh8I9WyhXIXNYd0nGGZr6rcDmkHZsl0RMjM91cDjs95ed4idonnJQfumK33FJ41CsjMVDOKHB
CqPD1mLQV7Qor3+2thpndRh/RCEP6O9hBWXkIWbi06OwZjT0BuJCDduov+w64sqXC5c6v1a4TQEI
cGluMcI5c2K8b/Al44hlRAHQcM8ROXnuC5NEu4UcvKUV8IgniPwiQ3eYfih7uQzT+CA8JeosSJ4B
KvllU5s64KoArTlaZlVOE3GQqmtkPOKWW85taCbLza0DvOyqEg4DvJdDKV/8+rzCMCjXe/U825k9
XcOgmmxYh7cKGTDnNxJ5r69jVVFNQP6aYxLAyo5pzflHzlxHNseBJziWJO0SHkTz+s8qX9Muwj2f
l4eWE1o2NEeLglAl0KF0Fjhyy9y7d/P/boHtH8MjlVf4obkKA3K6USZcvtRJ0NKSZL9hqgB9U+XX
ndIv5PDTnv0dRDsDh4noMgr1syFIsRzYqNGyoVWNqgnApuTbMYZ30h09+k5bnIZQTy7LfBT1KU1g
WDi+MGo2Wo9c2IoFWeYYLyBF+K3QarpyzH6Ba7OSbUdd5TfYEnpQmaIY7HrlKm22z8epF+7A2A8u
eDjiIr5784tQEizx1IP1i3QBzn39jF4OdjzLcIwE6YZWnI21nx6usB5fZ8o4aW+sFoJyhKj8Eyl3
4Y6mD7RAY9NOEC4soVw4R6/KpbDU5W94ntMHmzSfPAeva0ZK9ThIHgrULkkacq+1cuVeruVqOMnX
6QMk3niuVhJ+8zdz+96NpGkjzvOpSQQXaLH6nzRDLhvC1wRToVWT6ax9I+5EdxLoKX2y2vuPJIL9
ah+x1RSlzbz4Kis+n0nhA0S09ISWzyWXxXOerTDyXH2Zoa8jHEW/vQ4ZbthB5OgXdzaNHWFA1CT/
Irb0egspBRRHdNafbd8tpJ9CqocM7eOmj2gq5RLO2DPfmZzn0m/VlxymtDaBkDVj04HMXLAtzYyt
ULxpoR4sRE2D1dC8m6AM6QWa3OUT9u19r8ICWEFxVHpax2FW8ZrLT1lsIERTrlP2/0yNoMMrprvO
avA2rCp7ZMsaZSfM5hsd5J57DIukE7ULd8TxKxfglxCVa1AiE384NuogdcxT396nTKaGbpyXlu5o
iaTnAjbDsQHPIVPi+Gfg3+5edUNlurC6yoEjMZUQhQAqMgUsMw15Dox2dWZVSXQQVC/bbeVLf1ce
JmziNBtuyWmRlUN/xe+i3MPN0/RKmBQ8+x31ZsErsBf92ouxyEs7IhCJqJ4HMKjOXaufsAAqJI72
W90NFPHJRCV7xGxMmZc1KyVxJ6qG/oS5XdqrHsWFAsRbR7F7paYUPJBMW2lBnhfO28s4fQcRgr9C
PmfzGZR1b1aq7Nof7d1m/zPDBzM1LvIOe/HyEhjUcsvJtJaTJ0dU55wvXZIu7TsvB36FksgPdjLB
/BpfJteQUCYyz3S2DjPTrBG1F1LU260vZtoIn+UmyudN3Nf4+z9+PfiqB46w1SDrKbYNPaXeXzkQ
BIpn1irY+dIK+IrIKrCO3xCh7LcALxkLo9AlUN53sqBUFVjKLXi/0S26LGqFdnYimT+V9eP3RDwm
LPbZDLuZfZRsnUOWlVoVfZdrAy+QEb5rOlh8W7OfRgzuE7scNMBQJCTtttArEDhE+7CJ+mX9SnCh
pQqxxF1QVWDQafeMSVMKWnWc0lG4O7nRLvfgS5g9Mk/iSt0MAx6OMBVqzwirU9Qw9PeXvzvYZ/g+
oLBknpkmftKLysRc3h29PQbuNfaN6wRhoa/twK+24seXBjanpayoB9oHnBoN0C6fCcDKZ0JSRC1H
i9TtmjPmRx6IEkBnWie4tgy6sGRKohV0pTnarfYV8FLH+GhadvcBJNQUCjFpjbXJvf5f1oZU0wuV
Gt4/uUZSc2SVi9vQ/WIbafTi5x2xdv3FtDp81MNDtdZFT3aGjFogSt+XBMx8CeOAK7jBxiWrvhSq
MxMPxUxOfV++m0J0qhT9tOuBPWfiENaDuNYEkMGGJbUlj3l+tIwR8g91C/ItWb8hZn/8F1IxKQJO
tbMqSB5CkiXUJQThq/8YjvO6SyssmZiT08kRlwO9ANYMsrhSjXGauU+lld4TNRID5sEyZcTFsE1G
OjSfB+7V5lp2D26IhDuTQ/uDbqr5D4QEbkrkfUwqVl2rZ0WoEoMMu12AVtQ3ZPhtSEp4NZnsSr5n
k6ibWyPw8Mpzqx1hqnplrSrBSxiJpunztY3/Ra3Gea03aG3hHokrzqTnh0VXaygakDTPSqrihA80
To26mRe3dc67E/HU22dvWMC0FPA+6Fq2BzL9P+ZGZbx/8o6CHDrZtdaNpHOLjc0KaIg+6KKDAvsx
9ChcWikLq52X9Rdn1tfUSgFZM3ldBgPP6bvsURsgUOW7jtbeY79Ywlip0ZjCtMdfUF3P/uG/RHDy
XAxuKpBnjBvEj3zr1lqGlnlVsXhcotbSx7Ib87yo8K2jpxzbsqH4L7Xy28VAqrOCQsFH82+SquzJ
LHPVpzWoz24WJ3slDqHI0a1BZV8M+lr+sBLihRYurOa6fLQw00e68Jy7dX+HtoxhBySgi1tPHEl+
VGgHYPeh8nmNUnQ74LlX7iUSrwyvrEWTUjJGY3CFUEcMc1tPSUJ7VcPQd3BouXjM2L+Om/NDhoCS
ciFrlDKFRWpD+c7eDxy5KbVNy4QIAT59RBWTD88+5LBeS5nWLncnlrp9aBUjhthMxmvcTw8O6TC5
tx1GCaro0CudiLreI+9mQcJYQPCvsPEdBk8HAJ3x8zo8Zv/Jv1HD56Q+/vJFlIr+8mtmrfbEvkNA
ZZGno7DS9/aJOdy5l9DvuOUMQBn37Nbf3GQx1dx7CEG4OA6it8VeIGFesq+rzLH206SQb8nMHTil
VBj7j2yOAMRXjzCYGg5wJU7zpzKQwA25HWtSS0EX5iWdiibNR9UDYZ+mMYcDtRN0ds2GLLHlt52c
L6XZUq5FerARSXC+qvHUjKtrLvPY3LFlGgayaxL80oAbrisfEfPH2mKjs8OOZIBB5PtOgxH4Eo3j
0cr8G8Rm5D0JXz22ChsNwot0Wmq2RLmpcC8Ft7h76sm02Q1yCzyv8/X+kEeQr4+4i81M/cSuYUU0
+K45awL5JdoaYTlkYYUT7k5KMX1G+N55Z36M7Y7Sw7ViPmn8Fvntjnxreclxo/orqjZH7pNw6Fl2
180RjAxgGgi7ZABWIH0Rz/4dD4AQ6/tYEoPNyp93lcGN8hZImfQJ3c5lbuj08kgikSoZ/Oq0hnfb
eK9RiEfyDOtArc8QOohmTov7g76H+0Lq62t2SRwNuN9eUI/aM+N12tpA12ZAtRD8f9m8ZpPUVE/s
w0uo+34vth9Y/TRc2ySTaQt4nMgotPKyGp5Gr6iCRNGpybX8luAbKaP/OXzhEof0rSRtbXT/xG3G
Eeq1ImkiGS7Ou3qFe9Cs20mCXo+7I8mby+luNj7uUbMxPdio/jE0WvRFa53jR1FS+WgrFMTHcGZX
dNvYcIBRDoEHCqA04KoZB2EAZaQHC5wax0AbuXeLMsUV/zR2IKrNjYS9Nk+ZPnI837sOMU2wO2lD
esaUkGC60R4Su7bHMMv7EHQDnE3c/1mTPBQDwsK0nPuIG07lETSiojbNuDjiFhda/cAiPyfBhQP4
WDz5l2Bwaq6DvQhVgHEHdvriH0THvm04Pp5X7Ia2B+QZBJZ/uOiQRTFvCR7m2zth3JwWRfPtJ0rT
ivC6tLTbBBZ+9hlbUbIx6SLvJuZs3T+XJHlUnHcYPp2lfcooUFTxKD69yimj8gob7dCUHpeQ583V
jVmJAKfhm5mqMGZ3KNJCWtcTucjl8p+0ZthDuXbzkDc4bO2dlN7KGbAg4KbBliRFaVpa68yWo1AZ
Vr02rQcttlCLyhookxsLgyfU9QwyGh2I4KOj39qrKWuSHeEHnkZjTzT5/MsRN/aOQs0rWPiozNx/
S4GDf3Syb4vaMCZrLDUz/hcAdh6Eh0N0WxVeLfG+YsTrq1dwFBFmiHPvyKMQrm/dUbgnDO7n0GQ9
WWM5oFxKGhLcCx0nfdMvqHxkDDIttyVHZWyv/eN1eWaBjKZyks0ACRT2iRtA9wWiglrTpjOmWgyP
bSHwzwUNKDavblnQPLeR/0k8LDCWwtQ+E7rH2wRR3pxpEd9OFHJkpthhZKU6SPnszkB/4RGYzpT9
4AQl84lr9e0ckdNskN2pv+flEwpMdwKzF62KqiWtuitnstusf++FNpTa7RKGUA1Qvjv0R1bjl4QI
QPTdfufR2zfD1hdlY1x1Prm1hlpPfPkEIxl/y0E3vRbsVOJBX+HvSXxkhwl5/4IvowcZAYbA7Llk
nbdMLO2iohmFLLLjxHZh2w9yeJ6pvo/u8NHX65y8XH7ueVb49Q1U5hxgoafOb++F2l5fphctdLRp
VfuGQqNF2odDleLdcsCjWA1QQ/eRzQAIgXUmqOeu1Yck642VUcad2Hl7RZ34jG6nWXi6pqj0e2Gh
ScUS1I3di9Vs0ouKox4Ngp9vCTKUvN6MURj9rwvZkk4zGhPdiCHjsdVgYz4XOq0sHXNgyzMS5EPd
/s3Irpl/O8bgdphZCBhWcx6ffC6rFRZIW80WJPoExPsX2Xa7PVjHVc66yie2UbGF0QlLYIAVmBx3
iOX2wPgiblhyotUpCw3EB+jCmUFxRCmgXCKjTq8JDNIIvOAIuIQCFjj3ztrhheJ90pbkNaLLSbX8
P/mQoDcOTmMebgrkPJ9IBcE4fdF+Ey+u5bqWc4asXykt063EEDgUXNKigWKbPOk38zEGdPZqNw1S
8Kevm5tw9MxFDNQ8Yp6M0dNR6k5EccB9FEq5L7GaYBUUVnVma61Ee0GNgZt6vBIV4iM7qt7RmSgg
5LmF6WYxwjHRUhhj/T3mYKa3s4iyUPqd+lpiDwtS6QkOK0zyEfGtV1OAe7lgWOZsnK3wnZohkj7/
OqJ9CDCLNW0IP5RMiqcq1ZlArlR5ntNTfXmuiYL1GGV99qMBADFOE5MR5XahtD/oASPko6ivR+oh
1PXN9VqVDTHjuQbXt9+96SceXMXlLJyGjL2RbNk0mM6Vrh4inu09FSmGISlHzefgAkmUGZgUSE8R
c8aq7nlZqWMYMqkhaRlzVExHB+ih/NH4N18U0OAplZKKTZw2gZnEe79LFR12T+nzkHKJYRD8AxhJ
Bv5D/vao5Vee/n70LZtVsmJwPvKjJdssNSxhkEE4awq3vReUDQ0ul01oeIW4/NfvNiUjELYGmGSU
6KDiPOp9l+NEn8sNgEZGW34rSCZRCqnja7KftO4tWdunA5CERKloddPkidYRvCWhje1rFoSSrW6G
uelRr0bfUolgrkLAlnEC/HZVq6ea3QO1bt1fvrkYrXNfDkALCW55cT08I29+QdIXz93liJW9yAez
+KeaY/VaWIHiBhhpfOLX7Yh8tv4pSogjIVVljZJySNdOfIYilDQi6QkIM6OnQMbOZ0g5/a0oHbgB
xCrgeHBP3Odxj+FV6qzv2YuSFqhna5N41MZSxaV7S00Wb7vVtn60AKm6zE0HgX1hkoDU4REPvu/X
ApgvjZ4slXkjwqPkRxUJUKdLZJi94GmCbjVK8suvoe1ZVaiEQIXCPWp8jpDkgcztElNWdMuDCDPy
rMCu96VdxUzssXkwI0yIHjdUH4kesOhKXZFxhg/778090xv8dqNonXuZLJsCiTBMo8i0s/97K2IB
JNClDRNt7sbcAfzPzeRU1QypaCDsQ+vqTtlCt2SVIoibGWgduSU88wMpp3XJ23qiZa5IusrZf/7s
t6GdO7urXEzSIgsGhn6MwlSlUHrRJ2cRPo16FOVBw1ZciKBtz3ezyTRrBw4pZAwhsHfu1tWinGVH
T2eFYhE27VFVVd3Z9QC8+fuM5rnSZz+wFk2mJzRuekjenVsgMpnRK75n4RU9O3w+/GM9kRxZNYEb
2YtyAKrCTM6/wUm0f9wVDPTyI9TInZh+VKI8OvIbc7P8lsTyQ34mQ2TEgSsCH3MWbzugeTanngvq
PMOj4+m2x5XW2ciDGjAImhaoyd3l6HdhcFT6vM/w8+tabkVyFy3IOL2jlAY7N8aSmLny7zj+imrh
ZvS9SvRyy6YkXatjXlyxlrn8wQp9YNzXRY0VXpRH/tP90/4OuNTlw+Rld2oTXhnKouEpuPm2Jkx4
szn2ADEILtJy3i85ZLYzg8/m/XReB9GyNhZ66eIZjGQBtwUwjeRuSCFLRwPZ5KxjSgulJ4WMs8iG
Ei4+afLmp5CO0vTQqFxit0DnxJHxWvnka2y7aGu4tfjy/Lhl2L2Kegm+cObEi24QlsGWGJXSu5LF
/98MMdR5E3mwwaTRKEsSN4LB5v+UnY6qVZRJsVJq67NuapCytB6eQrn+sBPqPPWzAPh3Z6krPVhF
S6bMSrmmQf/38j5sFQnGDtZSPM1jD4U5GuddXskW4O4zk36MwIODz+XcQQLu/+NfByeWcle11vw7
FBydmFV3qmESstjDsqNhJR38GwJSwYPB/FyICd0w6tMNDeeqbjB8qRodxV97XpMYMXHu3RNbfMpQ
GEaTB9UBlGUyTFlVQwHLRvKGfIEUgOb3HYFVhc5R0bringXA5uFr8tQzbjGB+JpcAW2L4jYs/+nM
n6dF13gM7hAVtbOcGTHWNNO5xsFfahILJOoSFy3s0YwkahWySzheaEhybxWCUc5pDQD+cMhHQXkB
f+Bf1C3NzSPZ1ydfWbQ/eyODorwawrCfVXr7UdMOZ1i0wIPOqnv13g1Pl7eQjwVO345SYQEDJyU4
rT82OyM2hzIlxBangx5+G+mFzczcth+5NDPG4KYw2h1Vk7VDD8Tn12QvjQVyUBvse6tXELxKbq8G
aAUcNbCWis4T6/2gbh7NBnEkOcKCuF0LLE4WWioG9HFhM8AIXN5mbllHTUTTQhHgyPaXFMPDMITQ
AUHqC9kxDppJe/Yo24QtWPTG/ZilUv+EWkhCJ6qZMdLsltwBPY1gsd70AkOQqC+9Gb0WOxpaBRQg
NztlKl8/jQ7IDzWx2mrQNJf8TJ3Ev7viRAidVv1UopPdN5jgoM72X5dvbz++Od7Cx7qJjst70uIE
3rM5q0AVJ5fm6fU53ALhkL1//7qpJuClPwHwznwsUOlrA1G0an6CF2RQrgwxUlT3k9wD+4He9wqO
ilMUaP58T/1EVhYt6oAh0YL+LgGbZ+iSeha/OUKoMWcFGTY02iNtZ0rqadEZ+L6zGdhpseyocpXL
tNzqweZD/ulWv4+gZmL9RfurIBvMt1WyQmeCLwbTf64WvlNlgko/W7zm0cVcC6+C5/3FDAsfGGdH
v89Adg6KFUMLyZPAvdZ5zXGhzv5Qpo4a5QZo89g04SAnc5eCsix5ewAYh5jhp1CX9vtnzJFKh2MH
qBhBzde5tMyzk58drbs2JxU8OMfnEU8iYHQOSs900uVssbMC5mkZFn1eyv+PkEDl0v08hH8xsCP6
RWJ55vAyEuMrYoM15sSKeT6MxTRFBB0BitbA4ATFo0zwn1CuD+gHjuFp7KJ3WUdk6zEZqzBcHiUw
MmFmin4UrxhWVC3eKw7ak2fRlnaTAjiD07tO0UsCjb+ITYxLwSx+1Z0kBVQNulYoVxgf7w3P2R36
CGG2nOf2WerZSYYghV4chUMg93+XUv1n937nLp9vjjVG7JFUe2msbimzjHGvz9Hb37h9blnCF4Eq
RdsoJ+JOLe9A6NJaTOg5uXYAdbGh3Q/hV6r8e8voVi0mw7+EAFGdZ0u1tbA8Xkb4gOfCtKDKLDH6
SUZiF9EE7MLxmG313zgkxv6QCHGo2zLkbDeB0QIM4cPc86iFKUnqTl9vlXd74KWT1bQvu6+8o2d5
w8OeZ2HB6wWO9qN/afkrDv24bkgIFzQw+feu2+uqp6gHvW+h0PEvDsOblnZwA1BILDnbA6dAHf+m
KhfIdjiR5AlHg6NcXlKOv8xDKYrMQ9XloNDSHUQcLZRmfVLu/zJ7GSY0j1JfQ6OJ9ZmvSVdIMuVR
gAxSmJJH1v+JsfdHt/o3MIhAJeXyRwoZTdbXCaIPdH4n8vpTq4wFPaufQyCIpFDVQ4JURq1vFoMt
TOa1fZ0igz97W3OWJvVz7F+oiiJtUVksTVIMAhBTjWB32NyUbStLFTRbmAOsAHA83Om0TVKN5q1E
q4Du60L+/882G5Ud4wAQau1bPepSIf7MxQbuZv68ghZ3cH85ppESFWAHmOP1sSNKkNVBVNVoAOYK
qxwWxw4noY1t5P/Z+Irnm/kLWQmo0y8s6H+ekXn8Fa9H80ghv0EC00XiGErYItKGb9kYhb3F2kWg
bNpoJMeU99WmyJAPaWljOy0YoISY2ZcckMLzx7V/hPQATchDTYapCyIpH8eD1Rc+Ji3/CopxfX3i
y0dOyrHcSU7RsChmc9sJxuSFr5B2/mk/zYDGdY0nST33oxnxuhap343er3Q4m+PXSu2zr6FrEaSX
YmE50bZNqbwbebyZkpROecidTc3b5/oTAzhdO0Yz3Fj8UPI9Q5gBh3ilbB715dx5UsLG6dBHAzF9
xIyHC7iMCLvjw25h1ar5Cy9aY3wpyVLRZ1HpNC3tp2zPEFNBIrdqSEDfpPosbjhFmW6Pxa48Tox4
mfR2+pbbTyCVGg54fZ4aOw2jhiB1nGkeb+/v0SWQlgLI4rRcDLeV3unKoXB9zZ3ScXSTGVFIMjUe
lKLmZVCY2eZKsRJkgKakS2x3nslXnyCi3xbxVVSb+V8yLZpwsXTuL0TIIwmFi7kR8v45hOg0VKoU
BI4ebkGhDmWG6mzz4+E6Mbi3cJFnUz005BGEPB2stODOG7Z2wKApVglGcH30w3+k7AYEVhSqJfr1
oI36GbEUArRNzvoc4gAZepkluOjejBhizbW1W8/+GFUZfUkWmWkoq6OICjo3dWrwpUdv0ul9TLzV
w36dldmXu7RBVf3R8j+DqVWw6AZTsYjSjbS/BJrtautiP004W0sMCyx4TQ+fG6xPlE2fKP1uYONz
PHlbPZ1bPceQFFqRlImnaLIO6SfoefmjfbMsFuNtOSP63L50IbSl0v4JOGGYHWLZhO/OFRdDaX5j
ahNgWnf+Voh3g/ZW2m8ESKe+wbzOC0ce2j+mxYxQ9Vt03aADqOU5WTZG2EwujpGPkAc3MYrIkvzq
BTSSyC/jUVTvkOg4IP7oaUfgADLnkxjrjGyFrQq5xC/R5orVRYytXm+y2pHuFV2i8XV9XydQXH/K
FYRuRHdLcIblEQk7vs6/rGzMAMrDWOTPCxLaiA2yA5t5O8rYaPVExZCfzUApy70mACMVbfEI6439
+9rwlnHx0lt93PSLE1RpCgZl8waquVIrWM+JteoJcw0/bBOz1XUbfmCp1n9iuzwqYQcQMpHfN9zT
D4BdLkAl+Wxo30+Q7KLX4lf7OnKCXfbdgz/1XWoHzMKjymBvkL+zwWB3px9pWykhZTGw+uesKAv3
u4SMmMh18UybrFu7jK6MVul/40LEreBtKbKaYNHnFuHgnQgrsoCYceZOhPZq/tviuAJO/LWqoJsb
7Wb3L2RXunmXqCo147KH1fEsWjcUH03ih9xAuA4/Yt0x4VcC5E3SJ59ur6m2K4ANUz8wcqjL5rPu
WsKVRCZkMtaYXrywxOtypYBVqezehhHixdSyUDwMreFPWv9uhq1GuxWg47Z2vR4QG939a2XHwQxP
typD+TQjSMUiBL49thVfaoPzerIRBWefYABtIL9naXfUJimSefzTSgFkSQzSA5/xlPgiSU52/fYw
aDmuEQKXb5Gvim5S/OqsX9Mpkq+CQIyU6uHHIeavUz6jbOQyychRhdSWDE+UQCbDKm3LvRyMWVZg
t1xuQLDMRnooZYnVBT0RoCLeCQ9KR3NZb+CZaUO4Nm3J8NNieQZ7kxln1Mrsa5Ox6pdTu/IiU1qv
j6mv2riLlGng4aloguQmoSMHbrP4aXUEPHGQ3SkN2ZqadDOtWFHDJke+pbd3g3c6B1kDVGOlR9KL
2oAyusTRAxXgFIZZoMYcEJ/jUuXl86KF5HHNzQITghBMDOBuKwAmcNQlw4GxVZ7hl5rBhitkC4pS
8wvYWwtfJ7skxcIyc7QjPmVg/pbHQIyMgTQUn1t9pG38RgQ7Xjqgj8ci30ufsmk1Bp2Lx+ZcrQqH
MiDl9KrOFtVzGzIkpCxjo/a7y42uEllyo2atYUfjOXDz6I+3t7NLLQOa8clkUj6i5JQCiHVg05ht
eddpRtpLaRiGlAHjbgqs0jDRdVnmGh4Fnas0oQukO8XEXvgPXj5YOOhUSVwmbmpIXflBafBuYuD8
l5s2r9cFfSLzWDE1tQr/wvXt8FPxSgLWR1lGiEZFF77VtEsD3WM08MOL2YxgLQJ58jLD+QHGryym
sGY975a6p6bymMivHMcSzwN+qaG4C3U8tBKf2AwGj2T0fN+yay/pmpSZvB0m88XssowFWNKov4so
+5KhNQnAik/WO+cG66687+s3GpOmrcmYhf/164xZFG7QsOOcXR5sXF281tt/+mppPcC8mYaIKEl3
nlFWIxL0mh4oGJKQ5wpfP5uZmgU2C78SOY/oCNaQcxl7jmXflmAT14YYzDOtntfitXPQUbTdEVy9
4f69emntM24ulFVbaXPCwqTR5snyKgL91hcjDpbt81PjTrEDuN6IAbw/T760bbczAZqy2pD1f1W9
TAf/2g4J/vt/fyGssdJUwjn5vHVFWMweULOp1lawZ6djXqIZX00vpzLZcWKeBJ9wT6M7hqNUatvZ
VHunvgY8VDF9JC8tOEa662hacxT74H22/wadAymT/zkNuSRmz6wHTo8zMuYxhPog12Ngel6awjPl
Y/aHs/z0q97N3lUoJWbTvtUKzegtyK326i2FSm3BNkopD/oexBk9jeok53cFfNYWQ7fdN9o1REjg
zHFjUYUqRCb8yQoWIqw9hyNWxPo5OlFs83CBeNVZbkg6Kg9d/AkqOwbmQahi9xmVa4MOBdSijSCm
EDkeBOSsd3JXBUr2l3AQG5tjAumASe+h5GrhIyXqjF/fqrvUCrOcpCQCY5oI/ISeMVmmiStTvB0l
QYzUcyPAgD9cAhtOkDj3LHIsQgiS10p6gY8mM4WARfT+ajHUKWw6N2xzTqXdJt3jBneTxsL9/XeF
WTew6E0LGT+Sbi8+KyJTIHls5Rq192vCjoqqiSWETanskA8hJYj/SPLv7qbOxxofXFsVpWhnM/BX
JxgmL00rHdwP8kcXqPmLM7gv36fgJ9LaaZltRj7WlnqJTqCzQigjfXrXZ6lgiE0P8bUwsu+5nvDS
cp9iDPueS9DzyRhzJk7mkoBf1njI2gteSITkEx0tLqgkaaOXvEhX7ibcB1fgQHpFqHoaMbWVVQIM
zkiKh6BcLWRXSBqvPpyc7s1b9WgcIqC5L/AHcj57u3TkJVhCIIZWVSouKED/WrwA4S4s3p7mXMyk
ld5SIsFWSkQ45TcATjJhMOgMbUsVdKVkVBWUVOW/e7p9/QTkf6uJmA8JzsgIQyooCafKLgpj2FgF
yjWfWYTXtMkYbD4RiZHPFGuArZbTIr+N3gaNN7fsa4se9SAB/rHU8JbrG1ttchtSUdT2lmdkY6xB
S1kLHbaCR6Ppsf1WYWVNgYgdobd89rTWUYpA1C3UnDNb1TcoEladP54JTf9+D0F3aHHqnuPWcRXK
fz08AMgjD4D1m386XIqb4AnnIij1EQl99lOAEE+5yw1M5rP0/pZx4+A2Bh9SLKJAlu7MWDuJL3Tu
Z5iGMG0p3ZyGKJP+ols1sqKem2T/SfxDJlHrc4BVxNTqTP+bATDsDFBOrz3mtuCrMv/FOY1UCbbv
9Rnb8wic1BEualDj5YLEBo5lQmwwMuS2C10XAJNgtxEHA3XBCjtY+1hkyaaLu+SX0y50odRZ4V9K
VdDg7aMGzS6R4hGTtTPw1xCYoeLrPVFKFTaG4KmeJwByEivpS+U7hi8cr5eKFuJP6MzBt4CDvRaY
Zj9mWGXENlcWJJkZ7wMkBt/SR7zTGtA9M+hnPkZW4EutWAtVtAbJGBoh0hgYcBWG9+QO7Un2YW1d
xDAOj1uZ1lAYQHMZ/Wz1DJJSE5RbV5ukjSXdiluLGSgSoZdX0m4t17NXHLZkE6jLjuoDbQ/TEUwg
hgkO9zuFPi3KVghc3UksnZu3B81YJcTaPtPswPY6vul8QL7uBAEHMgr6U2GtrVTm3KiK424efyso
d7zAp5NoQaT6io0DOmrFvYybY4a5gujxh9kRPENj5jLI916LGNkQD4fah269qQ9CuBxSltwzYePQ
MbqZiM3iC5Gc55eTQoz4n5GJoY07vLsj9FP1WaksxdtwWFcEJHuUcZRMsiU2F/H0tmPVy7zCFBhC
AtY8fboAtBItcxm+BS7q0O7vSu/FChQM/d0BOaMgpJeScGunaZWLwXH7oRaBX09Ac7QEWfzYNEKf
0IQ3J67+fyylQJng4QIwuIeOSoAOWVhYaRaKRPqqH7iPr7W6lzZPyV07oTPylDLjXTOjke506f0Z
tWKJ+seDos0yEpC0j/PQM0rJuSyLiduA+uqYiOyy37QclLEwFaSrla0u1u0NwfdQegYiZlouuX/X
gak+iFZ1a4vm2siVis6KzzfCfw2Lh1U7XpscT9c3JMoVISwnJ9wWC1pm5RodMx4LhvIhRGaCcXve
vLfgsiRua1+EwNu1p1oilWsupKqO0X+IpLtSJqEDd25CAz+0cXPYliId2NS1txjbyq0sg91SPppp
00MLuPWzCtpWCGW8M/gRVTXSuLaDdzbi6srlcHwSqq64jZV5/w/TEZUbIO0FQy9mS6PVuSbBrYws
uPI8owKNAxggiAym8A4GKBrgI5hpzTzQCSw9aSGD9ZkMt6eJp+BVhJ2IyAbItcxlfIiIA+hGXWv6
h0ZE6s2kMTrS111KTD6zVCARbGcUydODqjBGhA8l03qL0Imead+3SZTug/WxhoRNkjY8IJxlRH21
KwJJk1jwZiRG8ODzDneb4dAXFqqZN2rZX9fRz9GVJtuEx0/23mplEgT7WL/4p26eOtBWZCmv1+VL
ZVjHTqoMFdvddd2zqqNghvdEn0Uy9oQa34LS7fEh4FoWbugkIhZvlPHYsR/wT8V+KYHJDBvJeY/Y
4ifWEIH6MN6N3PtTCaxsvsQHWkwebCatpvbLD8R4BDueFMgT6xHGp3tHOqTf2RmujnX4BC+wcHep
53ocxdzRfvYN3UChO+aTInPj92SWxzPDo55kaJ/iTV8j1ADHScc8PoEz7ivoMRmpFGtDrwS3xo44
5Oiy/8BOKTgwvI88GkPPhbtN54NlAH1MwBIwnqF12VS/afqmAXQcRtciQhQhg24twJakGKu/jLDI
R5kOMs3lPvpDgKsMgYv4yLglCSM6SgMFGJ/cULF7KJ7ZlIZGEeHQ182yGFC8feak8gAuQSPv74xW
O4Vq3qcghqigQroJrRJMGKMYUfQD8Xk1K6fo8mQzfZ6uG5P4e4bBkHdbnGIBVbd9hKlWTyUvyL05
tKj6uZXSEgnl1uaxuV9KssWhzU6V/b1pLAPn1Gm+IsTVuBzrTSe0JFxvFhUFAcveLx2HXUHsnKGE
Xw59BBdyy0s6V5eTt3/zRev8eJ+bMbNxRbZhKXjujGSjjT+HaJQXWPf4vgAiOG4O1H7PHe0/lzAi
6nFtugAQxVQaXoUk08mFGK7RhdLcr31+wf3UCdNJjn6ziLsFHdOYJWjZ0AkrqZd8KYJ6JAeKh//H
JjMyRSIiKNHnQj76uSmTILsSz5ZyKC+3b9DVXJrd644WSmyQDDCkSau7m1b2OW4MOgC5FkjVpDKy
TrmTTbYauSuPWUDLdpQu+A1PBZfpABjUs1mielEm6t6Qz1EkTbVqsqMk1YCgj7hbeMjgoeUKc/dr
Es1HDvPm/3+VvsZhGCKY3VlVQFmINMSuGQ41rBCTgZLfrpXPn+bN+BP2S/l98zrZTCRG6UI5OqBm
o19Wt5Lu2wvhCcAbAqkDr1p1sHZAla0lG1S6yz9oUXDIIPZ/2tWAXcGXl99r/D0fIVbwQL6ZWNqo
MvEKa862TGVFPSD1sHSjA/yG5rE6DACSmLWH7SyqLz6VxGyqEivrzcMOg61l3LpvxUOs2jKfgk6w
p5DKgOQM9YL8OeyM0NfY438OK8mXfqec7k5KSuWqbrgZP9qOTjKnC4LM3zlu1L3YD2PoQkh6T+uO
quHpYf2QtroRB9jGernD4E0CG93FEENBsUN+wdjzZD6PGduPPzSOpxq/hksd8+ZUGBzwqFFEPQGT
OAm2G6+d4ATD/kd40PSgV7EsBnkRWqWZWOxmwfDqIuQmslX2zfJ/moy5ejxpPMIDQ995KNPkeYGe
J3HJUYbJkKicCQB5soZikLWZz6V6wJ9vqjvqk4l/fhn1DHJ9We9z6B8axwkN+X+kAiJT0V3UXy7n
WMJhMQSBrL9+M9dMFEJXTddF8bcQuD3IW//DIw2K8L46bHX0SnGMttbtwJelMHhLVs4jhlRsKagY
DjDR7KBuysY6eMNGYaCZ/xvKOpj4/FW8xt3U+gfraNnyFxMgnfcfnQrxc3T5t89FvZV5sOVBvzPd
b9x8Px/05ddQgzBFR3WsJOcu3HLwxS5brRdU6mH3O1V1ggc1kSGyuP74EsFJCCNZUB5Mn9sl6G03
LfRsS4amSj6OB9D1YAnTkFpux6tZNKqHmmJx5PmxMA9p/32HsT93RQsdT6lL9zNNo+HvWmKlLECd
TgSkrznpproQPUyMVoL4PfbpCRCvj2jEJyZHEbgZuuGAbyLIAxF3laRzwTfwASegLQGtRI4qVYxg
ZU4NnvgT0pqhDsUlMVx/Obp0oBTFCQmP9WeYZHPa1WzF7Cm/4NIth1ZQqOiZca88Ua7w2kP3wVK2
oAZvFgO16PrrVfpzPwCwSZ07qhNEGZjJudsnfmUPt6AswkGr4+RBjdjwC68FEJqiO0XJvhNytb/K
UYfb6221Vio/IAb/okmxTfDhGzTo4C6TIRQbQsXSZMlWAIJufQe7cemliAYAK29PDhokI+C2S2Ui
n0rogcYNPDPCnqbbrh+F/ahKu7012cvD6ZyOM49gSc+HPNj1NvgRLe55IZIFh/jO6MWoCDouY0eC
EIolBM7PiG7M2+kHJcts2XI2tnjmshqtbC0Rs0olJZwpBvDD/wg7qfRCDjaZEl4eewUhaglsVr9E
dSdLNpmMvuJVUWmoZvmPzg4HqMhysA8itUphFoNlBMHQsri2Tl65oC1ZiBAetoQq4X36l+6l+WgH
wdSNcNQEc38b17u/4KRB3HWgu1e8S2vYpzBIHYzdQ3z5ZG//kvbQYZFRVzbHn8pD5vhTSz1huPwA
F9iiiWuUw9GErczvNgaMoXPqIalh68/14HoRxNiwMFSfYbO/KZrT2TICkGlhyq3SPMNZkfh+KWuA
ePO6VNoMzonmTQhrPw35gle8SzlrWzO3qrDtf5eUQXH65jSUoLs314/wMhFtsMkz8pkGCwBICoKU
7kxG7XdQZR9r2l6OXS87Ws9F9Cn1CnFULrYJGn4z8owr8WSV9JxSbgEBPu+Pi5Hyss+ctHLIE1u6
kv77UM62KzDguyQMmPOykOQzJ2vgQ88piU+TNN5cdQsP+m171QMnOWN95qVzoWUROdEUJ7skjsBB
lgnUU9HuYFVrv71bx3YQmNKy2TAWgBDBbQ7Dd/diVKlbiOVYQB5486iuMkHlpMLUBUpE9xAN9jgC
/LDo6hoH7mInwa2sSeRXJ/S1Nh2ywY71mAnUYxP+xVPKPtVPvkCm4P8ZkUp+hw0tvkvUQ+0LNmMU
02KorBXz76o/EJaDRnVEdEZrcHGfSs7UE7oQ6h1nAJJWfvEBHJN+GtWXDBaTwl+Bz+3REFjOuyGf
XQlWpdpyHSD4cysI7hR8+OGWSISi+1TvvroN0S+q9ZL4ubIT5FqdJg2eJ5v+uOR+nus57todUBew
JwgL8JwJlrOa2B5aXqNuUsUe2TTCfr0t1K00swbxO3jqXjQU/ukAcEYZsHd4XXr34YlVGGapoGve
T4nSHEfuOPf+7+ld5ocQRl4GjkNKVuljjL7OsV7TrQLZIgz/Y+uwfeH2BE++nNQC8GS1q58TjHx0
m0B1ZUNkjymr2nmvNjqO2rjCB3bA+zVi7YUBJYkAMjhTB35lFLiQ6nA76ss/U98jEki5VhVDMyUh
MJ/M+PJHIJ3YqDSS/KYFSySGs5ldQBI6pqiTUoT/xOXDlb3F8dTlxeYP4r5FO6FwRpHwHGsLxKFQ
+YwwKgmh+pjQx89nwYiqaxBaGl0eG51TxRBFImkHJrSNCy6CoM+qY78pYxHC7QQhBY6Y85OiqN87
OCiAnmsogS3Xr0jo8qpTL2H6yD8Jq7G0wsbEwuiuWt8lq3CiV/k9+kzh1w+LiLGCriAjZurhdtQw
03wXrHa8FYt9ox4Z6/+E1IT1fWApHKE8PYNA7EjzlFet/MLyMa9WzmJVvqGZ5IGthQ1Sz7vbvwJF
vwrDsevJaCb8u3+duL5o4Tg5j4Bk6cc8FAavYhYqhaRETpW709+OHJgGEZJGhp/9gnueh3UUs1xd
WXN7bEOpGyIvHNTPsFASgm6P2JozBpjK/2fxsew8B8Ky8shSbz/cFABpfggHyuVKjiG6pjG0uVcW
rcL1P4PvG8Eo32p/zqia75+Tm2XOXZtTgnXJKnjN7EtdQWLBuFZdbDx72Icmoy4Y5VPBTChhcoQP
XQXYlj/OReQi0/0YYCtSa/pMgoe8phFgQzYVKOL2b8q+29JKhaTpgjOmEfH7rqBOjSuC9ioZi7+B
TFE8h5bk5i4wuGjrLdF4LRrwbcQbraDaVPMIe5mkh5XFYADWfutanptsngF8eYo4gxfIqYma/0b0
Z4F0yiSu94ul+B2DXG8nRO4uEW5LnPrfzfYp7pzaB2wOH4fqsM6BF/wtOCWBL7HERe98IyTH0QH9
nnS7k0diK3vIv8w5XxH9nViL1ZmIMEW3/XI+fn9+ZRjYcnwvGY41Yf4EKVMbyDk7s40VCh7a5/VW
VHSY6inq80StVEEtBP6CP7xBU2oCuWkYajQClTq8Dmr3OaVfKcyoGcbaCDHHW+F95yxmr3QszEF1
EqfW8DpWZoLcUHeH7N8fcmbjVDzfOzknimunV5XpvfdB7GEviJHeitG1JikW0HhygdtcIcHYcofE
Jmz3Yzs4e9XXTnIB3W4b0E41L5ueumbflAj8gWFTSc0Ko7RPJwmFrmCY1Gml2ITtDlmKGoJC7vEV
aR7+4oAJl1h2lifhCAfe8aFewgNqod4QUS/S/3Wu4DOk7xzuQqfgbzr+K6vLgpJvJG4avZPhBo1q
AdBXSyRfp6uEE1eOrmAYMv1ozbEXZINmgOC+UQnLSCUSGy6cNapg+vduB0eLr5QWgLG14tM5VHSG
I5XJXOBpca1mwCVzarVyyBds8HmcgWStKKvcq/STvIO50C/1BtmYqUrGTeEZ1anpvNQVklho+cKD
BRg/pC6RqQy6UlDKYueaYuRjTn+C8bMx6n7g1g3tHFrhfBd5fX7ZyHjGrfgY4DVsRFkxgSd5FKov
iA4LtlVst+frzKg2nKJWQe4mtZ0TZbQBLQtdbTDASnQRsat7e9KP7miU0dR51uDf2j+NoUvG6qgV
8GthV/mSJNJAj4jcc1nGzdEeEnJI9k0EzmQwMyRJB7VIgjOb+O8hz76xQJ7tybkmOqhGa7H1wdbc
apLSPxWzvEZ6+fTJFVDxTOKSdxl0mMMWpsHj53xtu/hGf8FO0toxT7JjIh695Q1ninddu+12OrI9
iO6QWb2CetlS4651RJQgI7MG/VVctGHN4UIjLnhr1sPLZtiA8L9gxLYJLK3ZQkBrmrbyjyflPBvD
2e/ze0mBNNHhWm9hsfw66RKiZp8krlv7w54SaVnBiDcbfL7uO+RUFOfyzIOYcf3tA/WPxwWVMyOa
TrGvYenE68bGr3XO15Zo84i8bzGr/Vvn4NCWUyj7yl48PnJLVEaML+rkQHu/YSjLM+viZ4zSOthe
DTEOLnAl5WVPenxAgNuwUQxmhPh81k0G6HDE17gJL7UxnlwDFilDvZ3N9+doEOQIJCT46R/iHmrx
dm6gIftm35jy2DCS5VLb9g2pFQapfwsdk05XQkW5cdGcAflFglp+TgtphqsqrqfWxdSyrBmq6Y/F
vHdplIFRsG3CLSd1W7I9scWkHjaPzkAknS71+scfOJqCXXjZtsX1cXj8DV2ap+Q/Lmg1NH2zFWRA
BTinEPHpuIUs6atwMt5RxIUg2QEveNDR42kldKdVVX9kCBXiAhcB95YJkhtKulHlZkV56hPjy+3I
J9jb58mMiObYsPdoQznmMctJEGJvP8Jj8PPAV6y6yMwctbv0NAXLdj5Dsakat3hgkeVV7oKOHgWd
SyQLMHgpwK9SQEAUDFwSGtQMX6myyUNB4Pu/Fah4r/NT4aQgBOmfuTGY9P2PMo1dJjSt1apEoePC
L+FJt1aY7qGyPkVPgL1F4h8/9NfAxKjU1ZNzzzf+P9Y/cnU3K4JOyan7nCTi1OI+y95zgAqlif30
hMap9HwsSnEj0sgrUnM6ieK5HfhcxTwnwurxg3RPXgigd2N3VqsKmVl2KGSSBFjuo3RQ9PGb9/X5
N13GALifHEUcck+s32Uo/kIwdcAslv3IThzD4VT12kkRkglWgW6kHcOWoX4XIQcZ29MpAB4PG7qf
wzpYxe1IA1Pb2+kAWlNzTASesu90MznQqkWmIu+2gi2rJY2Z7U/U/az6+ZcLNkLCoikE7arTTAbO
FEHLo+S+asix8CZnkwDe78hky7nGrYc/jEadULGT4mNE0Nu93+e1Th/317zdtX8VEJphL8OYuEau
MBdoDT0YFeV6prEv47rtCIbZbVYUmL9q+k76PBTbXRmLtrgGSiFJVyuPVNJfx6mhA+lFr3lBewmP
1KjSOKwwc8GeLODXAUpZswKs7s4XdsrF9vel3VB1d308XAKdsiI/Zh4hc9lYI/uH/jJUFb0Xt/qU
D1d0xLkpXsc+aXvBcKPt7GGSTTc09WAHPEGnul0W9+NLyKO9MyDTx/yKr/iO4DUWZGEydEAA8teJ
nOey8YpItYP3hh/5oTfWLFMDbERAEiqcfc1FXqp4CmcOblQSzints+iGVQ6SM9rdFym/RWtUFZ9U
+p6b+mOwckqRWUy0961Mhx0zgl2rBW6jmgZMvKXoaNgT+wZnAJP7QSOArtrM8rZBRBR6svwE5NAG
kZ/X8+/nQxMh380oBxaP0XIffTdRk3ddO1P7Ze9lkzqiBnFS0beM7xPcZ5Tch0u6WK0mfs0V0abo
0MfTXPWWbujc2Wl8MccH7+vCaezRgfItivPVjEzVXLFhUNUfhJQuzZ1DYS3dE+aRarrKOo4bNKpG
dlkmb/WmCEJfg67GnhZIDNJLfO80S282OY2FKJQLlj5xZBcXT41NvmrmHcSmwBzKcuMm1ENjSdyF
zqK0CcbeFjqvXxsOkYPHCB0AjGdbNmPIYuzcHDWOZ/e8L7urL4iE9q5s6CKk933i9I127hUvZHOY
vGC2R+LN2q8QeAXtt2Ophs0XB1RhA2BdprdiXf0i+2JPs2pEbIAbeYUFUL+NO6AhDCJjK0RoesAO
CodeQjEI0HtQ42ykanBG3qvD7eAWN6qIE8jImNJBp9+BTJIVT4cJyQvHhWWG6oITse+S7MOwDYc5
imp8R49R7cBOld63I0+ucbI5YhGGcZ+vaBwyGyG5vemP2FWo7B5zb4T/JEwVd1O0/l/Ek/F8fPRU
L+cFosDZoPl5jQSBxGzOH5norABqmdojO5cYh249EcRjKU+XG4nXq3vLrC5J23x6Pv9RBe9tp14L
yG6rvQoFEU3Z+A2Lcrizb+ZTmx+F8LYNb7WlCZN4Zx9wpnXqzdciuX0/PEoICtR+qfIb6kgoGthG
TwP/cWim8XOsiSfm4U/2+juQTBz3Q/REv6wRrfAnyG2IOupaBxbVnmDwgP5jrJe7cq22pAmVzXB3
eiMqyGiwDsdFivxmEthbAqvvqRszPy6R/qRB2wQmoLjNS44E7iTXgbE2l29RC5w/0h+F4U61DHYK
qlCVHdgwWmoNhvNeljucrgIXdeGAvvefCEYI8zAbbwE5inbyq6AwCkAW6GuO111jLZX7rKaEPbRa
W9sPOs9HXI1VB7MYGSVd8LwFmRLr5gWQ3UrJ+ddI43Jwx9YEYsj7kGeEHk2GHxwzy09FFlb9+xi9
eDz3mhJQtrOywD9GYx3dVG5kkaXa2J/13RpWAHSqtonJjJ0tuNcLEi2IIHiwL+G/LlLBH08DE5OY
g/bRLFtkVGIZW/Is3MCVRv+31PgX8msMh7p/qbIJMLcFSdhQDLR4ROd3+M6oG4f8NKOiwxFL3TK8
9gvu+ZmNfazRCOLZ9Tp85k2oxoGWrcAx/X+pr6DKbUft6No9zdffJq8R+wmvWqR8R3AnHCVBMDzK
5vDrL4EO/3Bo8XghxIIIa2bVMJILnK7LqqXPtpateZz/aXkG3tx5wRfoMKxZAKl/81scmjps2quE
Ok9ETFtLhQjAQvivdXRbT9AsNV7Qt5qTXB6fl4y0UmM1wbwfx3mJbkGhqzbeOvKJIe8btDXZv5Hz
fSkyum9+q35XJv1GHQ3VMl2j8JUIYei/jA2uhK1I+wZCZDlP4ZIzFVHg2GuO6KoVCCHbCSkLTx2w
p1UVsr46ggrVCy3QJgD2+l6vcPYHXYam7duSZEUUIaH/1T0WbAVwB6BFuTrmQ2829pQ03C+EHCTJ
0jJC5GKwkZOwL7LyAuUiuUECieUHHnilVMLablPLgD1gZEp1fYsdh2bdfC/GSBhQ/K1yK1B89fpT
gMAfl/vuktUOb3Z5sOJ3KX4UNneMJNpTDkK9WMTDpzPa4kId03UfUcLx2EyV01FG/PtWJJZGdzxS
u7cZ5cwwOSPUW4/VqBdXrq2rj/v1qkeZ9utLBWOTg8eC+ftSFm2sJDotoDyPokpVMs/W16GDys6b
E5vxyZN8ywPJdzMUMAngNu2dK+nNrwsS8Sy0mIzCVqpwXNUBf5fXiDuhvQVK9m3gMNWMgXA7YUDD
+8ueCcrE2bjfkYtcBn6AxWsASiwPc3YNxjp4pb+hhqBIMG2DDRsDTuIhs+7P8SUzUlFSeO+BLOcl
sB9vmXRlyM2R7Bjq/D6dgbIl3+0+OPi1rIhQ2UDqv2TOe9WPKanIHO+TfgPDwbHwF0KS8mOmg8Rs
S2MYFbVORLQHBxj2RSsqBWZfmSQ+LC8LIzxyp4aIR0zVY8TItjfebJjhUnqqSGckZUY5h2IKGuPT
wVJmr+qI+R+TXiwlF3CI1/+k5bD90gprPlJSSnK56kMoautg/kusQBISkQVM1mcjZq7DM7qZSJmZ
2PwZ3nl4FZ3SSa4e38k9mJ0nNhMpi2GzrhvYwXBtYZ5kREHxLocwCQ3JfUnjFrhBxibhmJ2Hdz5K
EuWXCrjJkyw6nbfLC98dwvKpbN5f59eGkEu/U2iZg4f6NT7AYoyL/Fg5m2cUUPKEAMyIV74Rxqxa
Tj+mGHJI+LgK8HZEh1WzHP0NHzeoMvpPx8kG9x/IwzMQKvbdrPphmBeqnle7gk3BHm2ruGCvAl8D
S7sYtT5opJHVUcS6Mirs2FmiAeFhu8nYMc+GNfsPCrkpecKDfbvDGdaERaC1rkCT56bTDc8xMWqy
BzQDJc2xc4poNRUzC7rI850ZNZw29eHEuAIRrsQniegWtoIx4+BKHBzcXGuruc3R5RSCYEErK1fP
3QPTPBLb8j+WzbgvABoPkx+afzjuxIcpm+7iyNWZt7Kwn7AHIAD7yyIHaxDV/I2Mb0gTJMRzgH6k
YVAKcgQbj0IUyST97JUsiyIgpo/3ncItmV3gIMEyL/lZaa2w12TcsMc8jyplq7oqzGicnZjeLuhr
T1BJoll+kemVE6jn/8BbadM7NcCEvYNhQ8eKF3vNUiNv8kaUsBOyf2vi6BXk6lRiMhyPHaYzOgzD
lWXtwbQPjdO9tkY1tqhYEF06yuC75p9oEctel16jyXP5H0yj6NUsZJNNngBvnNgkf4a3bHSF2+1s
cPKhRZOzWVXwtR3+wIdn0xVdjeZRE77gP/u8Vge0xJly7N8tGDXYyNYTEoV/naH5vg3SPhapNXrg
/YZ/m+jf9PfEIBUI1K0g7mgZoeZ8JO/FfHT7BhtyxwzfUnbrPvaqivjKo9+q5URc+bpv1XRfjAlT
9B+Z7XKzfUiNazlfBIWIiVuRNxovw4wuRp4C2l/GmypM7hZgL8lwBzniceknndXlLuFPbm8Z7AOp
q0wVGE6R+gzt9L1R5oB+6tFCPveqvBeO0aYjEzaE65Sca7R7q4XwbaD0fTc/3XyToVRTxtsis7nZ
J9mswU+c5xfdFVT09jBXJVOnJK68pa+gTTBZVJYnEtxV9IpEKcFlmn4+JcCBr1XRyDdm3L6Xtgsx
hG/2IRwF7EhUaNIrSQFGP5QNUr+M56BB1tRAd8h8+IQiiNal5C5Q8itSrOHPD7/GRgvITnXEG1i+
U0ztZZAJ50ccRr0u7Y43RFQyzsrgZ05W26Nhrvc69YeH9fR7UTWV0u/rJCLdOlYPt+0NsXKj2GMu
l2/QO1zeQs4+m7SqMcl2Dhmb8PKim1ZaeyRzLHvgb8bXz8IFWR4ONjPXbLujYWYkKH9MDvsL0eRc
Cy7piYTg7uKvjsMdBwNDZkjxEsN6RChxvaqQRRvhIrByEBjpNTbQqh13zcTLg4tmXibhz/hjexaI
ewQkuTDqJQnDmfbwmNvrlq+sSagVtBVC8gRwlORLhk13/WxcdmqOc3Ll3qQvRp7Qt0N116NApLcX
aXhnWFEIR4R2mrPEX8o0H4k9LVUMCdMi7JVE40pcS9bRZ/BUpmRcdQPopsGpLhWVyMB4dRl6rvzT
JGvSlwBrFwJgTBwKT4TQd2cBqKRMzlfyA6UFg5NIFPuGeuLrKfbxecr1qEghSjrctLMBHp8qbWX4
ojXj4TSsUFxaIjzUwyhhebXeUwOt43JzOzH9jC8o+GzMKuvhJHBJ0xQwZA2F/3pYPXLa0wevhbfA
B1/u3dEXqQjxDqgYKWfkXh0oeITIpFBT4/+cFba5zC9xvNnf/E5uxGxzB3GAnDCfkzXD6o9SHDEV
I6Icr2KzNeyx0bWNPvGOMFF6um16s+vp2ChCc1vZsq5GL/BoBTBGqhgyDq8f0sMaksj8c0M1G8yr
ZQ5vFgLL/O4n62qv+nLpvDbEq1yMoi9E/XXd44pSDeNn3WRy1oYsZ89VrwimoAPvERU1pfEMWcet
K/O6Y4ZBs6rDE5cLIgn+yhS5Pk65G0102hC1GTsa/egqmE95knoCuszNmV7an5/XwfnAv0V7f7n0
8k5dqiNl5U7+dAE+u1alNoD27emPQW/RVmaFmUqJ/EQV0JhTzqCgECFVWCSPA7ho4tpUUGRZV6AR
TXrfFAEBlu38X0l7NjbNNjaRtwvDxagNJ1Su1786WAGb44YYrqvJRWzbLVgW4s2KJsi4ZguXh4ez
caqkDC5SPvRFmyjfCmWeum/5x7m++xbPYvirR+iAlvLgXhCIPkqt2QEPbp0SlAOR65kdkvpZwvdj
3CVrCjxIN+Hiui5Vr1T/Fsk3mxwmeGcEvNKcfaqrsu9Gvvrc43E9dP822X6m8jxpHTsuNttxpar2
AlRc5ZUiarJa6U0DVp4hrYQjND51mGH+jGVJi66+OwTgYTM3fd2g4Waaj+DNjGpErakwAypyXE+6
5QOPLqV2v49xaJtHVkZ+4dqvMAezcIUF73JohU68fMyVZur6LVztiEfZi7vWbVPqzbzAsI+H++Nh
cgQDXa82JlxRQ0rO85emXcJdWG6x+IIz0SEX5nRp505icMEgxqdZ6Hulp8C6IknCZVSV9kLvJjmc
0lAwSR3ObzPt7fqNSOnViR0GhIEj8Fx/Uaaf3qDh3nGCcZpUW3RU1CGQFL3a7XP5EIWfTx6bn/gw
SyTypkWCtvmOJy5wadgKvSiX2v46TBoTM33imFUT7PFb5hlkgqjwL39QxQCp00+zd0bwFr/X01bp
8eEt4A5oEcInAU1MH+qjMapovGOY0zXeDikLDSSF7LJEBj8mZE7KZrdhdf6SbPE76PltAc9xGJjE
ilSEVY4gyhcBlJ62TnN0udt7LndviOU3KZAbx6cjWSakhQ2W9StxE2vvuQFc/fRKaC2AgDodDTMN
3reWsbJKm/VFn/AJb9G5+/VYC8rWbUyGAPxetBMWHISrEE2f/OoNUOFxTdUG2F0A2Ry8jjgIgrc4
0q7VWWgu0cpNHJZALCv2pcKa5IR0NQK9NQgiFCBaovUzPsrFRxujqdXr6AoPDZ4gbB9HTFFHAj41
1UA9fLpScEPP9uoUcN0dOIg3AHa9wG7T7y7eaVnaa5HMFTn1IknN9NTE9sxNfeLCmlgW7RciaQ7Z
FIieIyvYWlLyLiqtitD1BET6E2ZETQHtiewxFuGopssS4M+xQncdwfJfMANSDeZ674pjMnsCDfKB
VQ6HmuEmcZ5/9VzfwVNLIIV6vyokRaRbMcZPXgZcWXZUGcX9uXr1cEebl4Zwep3Y8MC5RYVgTZRW
v0OOEeyGZmXBEQgaiqvi9CiqrtPVRyl2bnK98jJS4YXZCG1Py1JWhy2Rjftj4XluVx99W2WHBtwZ
BXNFoojTCgogtRz9G40uql71d8gPpksEFkvLlFUfr0NA9RGl5HXZolNX+hf7deXMdYS30uFaqi86
nfe/x9rzbXqDUmpFlYpn2XHlgBMQHVOFLMYiNgCRQRHmzc2vvM2xe8M0TgsWM5LjNwOkWmpBydHP
gvh42lKPtzt9m4IZZY1GcbDSIqgkNCUl1TpTk4vH0w/Awwj2y2MkT0FD/HDCivx8WSCO6LX6KSAm
Qv9UGvQeVOfq/MAqe9aAxif2uofSNhBW3+w6CEtW7Ap+1G6xxzY+N6ohbOaGopnXHdL1CgY1PHem
qhjGwMxRUZQoZZA5TewV4T08KgOlmjLuy6swXUfIVzU4Vg5stw35nwz2K7ilsgOmmWviB+R2qxc5
Irr+KvijHrRedwqfjuQVnuAlf6Cry9/hC+3zSDK6wsItj2b7y0AN/82ySWKK5lAV/YvnRcFMqFPx
uQKoruEWoPaW+UXNdjHl3U0SOdUNKBcpNHrauz7y0iT/HmzEJOUEn5vqAgRo+trBkzkYl5gtmIlR
oLzaC602fFcAU3hZZmdGg6Sjm0+aS1wYItkWOPS41NZGtPaQKzLdyezAXfYqVQEptPGH6dKgg7cU
a5SvtUJvHWo9bRX9BijmveV+UUZ2HRobzLdEW00of8C+qZMMKCHwP2iv7GI9tS9ygeZvayDD6F+X
oBB4pVv2Zh7nKUbmZdKenGcrIZIgP69S5Mu6InzJIyxhr1P7w6PglzZL56v7M3xiEbQS1LmrQ/xt
I0gS/u8ei4++WR8gxHvrDcG2WSHBwiBq/mR2ZWhAmKh6PmvRafbrJGaTyVra2QD+uxRuROZNMixc
hMzy6cnVq7YLIhocgQkpqiSgcm1Wuwrr8We6iCgcAX89FwUePDDrbPjIyTupWyhwh2mNrW8vvZk0
4xaP7BxXyZDJkASuE2sUM5nTCTJeXhaCwgJlAxqZ9osUp5eItOfboVK0mNVxtqRVo6K4XQX/GAyS
BPGgR1owk1FT+gC77SdrSkjisSaZ/wvoNF3fEku9mjasMWOTc7Lg9/SkKTY5ZvpUZtlbVTjNvjZ6
Lt3DiRlgkySBOfAv8+ouysJ9mPOhel+4P463edNX5Drxj0VZE0kKXshAruYFHvDa3mHhFoKSYICV
EezuQ8xySlfKcT8d3KlhAXbHtgqs2F3WqgqfsFEKP1eOVQdzhjeYFf6+uKoC3oL0bakL5ZuRlVmB
5C29sSKHTrlcdv7oO9rjrC7P49nW0xbQERXLNtFQ+SYrPrhoEEUEghAIp0OTYnyCpRsb5AKcpIWX
nNe9ZVDCbNtaqYNuUBjVFMF14GKF/e4MYVO/BMl3i+iZ5QzLJ7m4cNgqyPybHvQsxkfMkudpcoQ3
7dCV1TDqcJh6VbPNXOjXTewnPFRYzzIsKaQ7h6wQ+aSr3pQJOXHAW8QyheYySqJoUf57TJfC+nbs
V4GPzg7+ytln8xvH61p1FxLQcwlI+F9a+feyYsMneLHH/8pcBu+moUpW0l+UzZkTs/SQ90wfDFnh
CgZl+BSH8h9dDm1Bf15Z2FWmqN54ehdvURqujD9NhltM9VPqJgkh7ES34P2+fdzZi9lNMSmuipy4
XGxblX/6/1+o2h62K+L1cBphK3ODWsQG7vhqwa8fsBWAc/xHbR4swUz7LjeqbsiItneryOgTH5oP
SLGj8OEO7pAQl3MqE8x3+pUbtXZGnROGnNsiHvdgBDX/UOs05VztuSq7V4yfcPK2rzraiqOCFKJR
9nb+jQVNNBkYV2ePkT9rxxLgN81prmnMwqJr9Ij5eE7N1az4QHmnIEa2bsOXkVv2v5ba1KuwRfO9
EIb4J1RWXCYN76TN/YlEJl1XBc2RbIqs57celEvpVpQfyxS2Id5+F7qkz6Ks2TLqjlQBLAAWED57
PGaWCA3gRVYVVMpxaQhM9SPc7FWVt+gpcmB3yNsUFiW2F633nZH3rnpLH/MPxlMQQK0bL1uH/YVJ
dDjXxackoAZlRzWKTw68AGU6FT6bbozuaRRmYnEMuUytwlzc2gLbxknt8Zqeh/FjDsbiuaD8CQq4
3+TxxuwbZWg8upvQPhJhkvyVbYiNhyLBUKI34cp8SmJUI9ODI47hun4n4dFhm7efZVBw0G1d6Y9r
K/Af3eATcVsnjlWoMF2ztSU5u897TVuFaO/0d0q4dKjjWNLQRCUGH+jLWcm5KM88i0ltS2pnc/a6
/fXyJz27oRq27OSBNgMcePD7cAbC74BrwM8ju3HKAgsp7HYBVh45Y4j84rFy9Do9K11xL6F7E6cN
VaxWuz4yEQkniZp25GtaINMLTweBo2JwDU13coRa5S3FvBICTB6N3adTWuFCVQYTpfkth7J0K5nu
4m0CF0O+Q/t5TkJQjnmKxdfTB2AkImFVBWm3C0KmoUWa0SWt4LfjLdloMWvsXrMkUSEA0i5dRa7j
LPz1DPv5U4JOs3asUYZHxbCYCNSOUpGgnABsBwgeI+NLMAChgDukb3A5fRcNmiC7h55xfn5SV/6+
GL1Vomb2xh10887FyhY6Z6uatYOvgwpmqC/DMOwsx9pqj5D+/T1dbICkKGWAhSfcJ/fqnLqwyu5r
+flV2YbjzzZhQIit5dxsud2E8MO6kyqRodtCwAghaZXhiPi+3EtN91RsPAwxFh3uFRqplPyKIY3H
8GflW8emBTCBan2N91UVMGQht6P1IXzRmDQ+h5jrKOstvGyKHJnIvtj4B0OaXgdYCjpo5ghFkmzm
NxPdk7opW+IHFvqLrk4leYPnjipaV9VGwLae/dbzy1utnMIaomY92Ax+LVzasanzW1mkYI33GndX
7im45A4PPNnchKTC9dWAfM3P48CvNOp0fE1feSCT3IZpEIyTyhOE4vjWkVLdZdNxql41SHcJh75v
YfMoXT/RxjySy8J1ShhmFeGJU6zRp9PjMhTS0pvdlSeMh3WAVXOesdlQzwCNgc7IcZVs7EO8WYkz
39zPqjDys1TNkDERl5RfqDJtXzqsbe3fkIaEaWqZEXcwQDZntST/W5HysAkgrl7Kd2g31HUO0Ys8
Ui67zlYp87/g8yBTPgydiN/pkiTwlqKFGLpE2XfJmXVIEozMNm9DPQO3+2D8WyoRZcpGPVX5wxl4
TQ9epsLKT8giJfOM3LoEwIGgqHySP5FO3SPaDE21gV+e0AuY8+ZDE7EQJDxkVg0KD9q/2v88RH/x
G64R4kPH7kZjaa2TYPKzA1K74jbtB9vGxfXF+Fd5nS82YIAgibaVUFZTSBHqqgy2zCO9IXXchv5Q
kbsHC65uJ42qvLkkpHf9cxS275VI42Bc5QUPpoY7TUG8AOiLc1y5ueo2at4gbubfLAeRBKoyPLKt
u6Toy/d52wv++4G6xng8hvgVYTGVuug2YVOWAKo4tKrIWmJOvSTlF2827KQvcssUW0MXtWYcJuBL
YL43g8n5tsHOYgOTUEYUY3uy/pTgIwPzVKuOxQlsn1kSjsKv+5ElYPwLCXq+zXc4pVzRKjt870Ns
5N2Fo2SN3KC0Vr9dDkOC/GwE3wDgAmWAswrdTa3dZ8LdTWd3P6/mx/fMLFxHBLKjQsJCERzL8HqY
HrOVSslI7OpAHJdhlnonJOMOts5DVtfEhoGqCJcKaeCeg0AqyCqwNtLP0ZAPfTBWNm+0WU37d9HY
+PjUehl1/jtVKtGvbkMyU6Ow8sM7ky39SUhaxtx+FvZ4z5C9S6ewJZ1v+FCwN1YhXfCtxX5zF07o
jbZg+3lFpTooJLrjCbHyJpuFpKAHUQErRFsSuRZFvvJN3yU1homPsGV5om/TfMPcV9zuHs3qsDx+
jydpocGYbpIa1ZcYNgQ6i3n5DBnJeVxr3vRK0rsK+Duy1GVeN16oiuClFzRzxVvMcWPa34waQbGI
/PB+SmIOxzsQRyTgZ5g1D4gI4lIiGdqyRjmLgAolJhiVvldIAL3mjm99xkf7drII/MGHGc0z2uCD
t0xQgRXzmGZiDd0Exh9pFhQsaud/xAZOnCCzbqkMuGXoivF10RrLjSw6jyugpR5WE9iNGpu0S1GJ
thUAOxNMpAiaaFqItvSYiQr/dFqkYskXYv1+/8Hp20q9TjZxbQpII81TNyoh/20tJ+iUpP/BFiDy
pPBXGnEplEu5EjjI3nG/TC0IIdJw/GNHj7Ai82v7vZBXjR33R3koKIoxmdpOeEr+Wv+6vfv97U6B
J+MunU/+VjtxfMaNKbK3qo5lwWJvOuLaYoYU4AgveBTzoQMQUR6L/7L5Y/usmGCqkx3XMe4PM/8e
GWLFXAuT9aVbM7w54EZu5hO5nPqP6X/AwDFfFMPCibCuCeSOBN1OTDaaEW7tGNP3i9DWXSSZY9dV
xCiQbDevFRM5m0YPIa3wLsK1M48XOTZqPtW+VsSVSLuFb9+LECji4RoRiJjt2UZqISQOTyoAK+DX
aXlwDUI25+8alTz7FXk0N6Cfhx7cymmL0Exe6zVjav1Z/429yhh/D9pWTaSirwBD3oHVuZDmXsT+
LIhTB0zWhr35hZKGw0pJH0gef29qCn6VzYU5hOzd48u12xlS67bKc+bsLzTZweb/z3ZBhkBqFdGm
1qbrAoVArrcBlQ93hzQ4QwHLCsut0RfazA5HYWG3OJwEndReDPInp9E5d2h4bHKkYhCLfcFC/8TH
hOIXDMdPsRylYp8BC2EeO+LsjXqMMa1U+n3FCLKzxv4+UBDDSkK8VdE5hKZ9oTVpjmsG42htSsJa
wDszJBk9f3RGG7E1rTSK2/7LrXkjr0FGrLGvtQQVEGJVUjiebD1FGfeSteBmkgqBkgoQh8xfSVOZ
1BVux4R+rdWrDYpvy0kFCsZ9emLG1tgr8uLMH2IVwKFY0H9HSiHk+byzp+83w04T2+2uYCqJWCsb
Kk3dY7dW8I3xWEVxK8Kw+5wTVjWxlImxj6RRMvdTtfpOTWAHfzpnt4/5BocJVsnQetNbUPK3UwH0
AWhGWucPZya8MeclosD58L9jT4LSqzYvBcvLlxRfokW6lYTR9v2laylDCHkmSwxSPPVPpCw1nI70
DBOS9OmkFg2q/s66UVIUQtb0Kzycuk6Y0j2d5o9wFO2WKq8LqkO9acHdjCSqt0Pa+Ef4jX1upL2z
wjw48gg3O4YoIkh229ui40+zD7JX/lh1DHqauk93BgrnM99L5jC+BdkE+2ASgiCHZJso9yzOz/cu
RDRH0RgFPIwdb7V2PCtqsdYweEeeOSdo13S7JXFNMhiDQCa+JgyNZKah7IY1aH9GaI10T7GEalXd
BvsGbBRpNy2zsf+rSDGVXdgeKHUt4KLNDm08AnJ1cfc/p6EwajGlBXs7M9bklCFbVjkUjv/HZjg/
ha6GAZTXj/XM7DNk0UmRgY/8YKOa1uuvghMkrtnv1sm6okuSnRkHX+Z47UelgiZXasFzchbogIq0
7U/OjgLPz/NXnoqabNQnZlTiukAl3dLTherIuDVDFI/Qq18GihgGxDpi5Y5trV/1euIlp3jM9W/h
+dnGRDn6gK1Dyz2wB8PQ+o8NbijoEVQt8IndeCNrCHoFcLRExWbCKUGm8abDujG/dG6oSJEh2/kY
oGU7dae87N9EQCmGrS08MxyDcWJRgHPjDG0VQiSXPcI/KulGLbcu+rpBo2N7qQD8I7yUJmOOFZIM
T1aMwsfN15GqaFpg2AeYKgBHVuLGxF5WBCQQbH1lvjQiYmctUPLoRcWsUD+aemzSbaptVCwm9wX4
P0Mpqr53SFsti+hz6ooy9ZP6hATnQwzD4vhiMbOqRS1guFgcXWQ20YzskAGwqM907qlR7NTgTB7e
7slGxMp6DEmc22vr9bgLpuRzQu2AuZYS/B+ptwbckFbXp5VTQUdgZnQjKqmspciPIYfpKPhU0vzb
GnN9Wd2Fb1KqLZpHkxmvc9vPVc6I0RyINsrpKm/DzQ9dRAs5zPb6om9bmspUKUHZx1KffGi6zrWY
wacG7IT5SBirCfrpIKPllTpoxCE0GXYoNRMxeTgzNOKWJODL0uVpltHwojYBreigHP0VeLw59gEX
srif1Iy1a4NAphzHdpL25IbAxhHTqcX1VCIAw5NJYJRxcJgm+zdgo3LvL0SI9eZIj197s0NPH++b
q1T+6DT9yHQs+IWTlkvhlgwqD6Qw2rwgEDXGGpIc24BDRL+srDjN2A0FxAlWfPVfKXdDxih00gER
8Hq7qBJ+JgTI2FDVAF21D68TtG3zEdcFpurT9/7LJF1F+o99aLpCo86lpGghBw3ezZY9gCI0dRFg
IXG5aeHEP1RwLf+4WXxRphsI4JXhiey/ZDiNerAgIQnpzsz3CKK1vAjFi7pIzdmNPeCeFqNU46nl
+01iiSasG+xJpTL/QU40NSZIFJV4hHIR/VQqhAvNiI1GuDWggHILGLTcbjZJ+HOFWHBXTuihcPCt
3dBW2EjZ85ddPiUZhRKqLFL7n50qUKfvqjBrU6f85hvrMARODuAAbAqqaQQMxTU61dY5EgwiWM48
muI6U0KHmrMcyOMaNGZ5RUOKu3LXWNAn4JOdZ+9QOnO5VXUuVDYDOJ8c4kw7VyW/eHML7YI+KRMC
rm2yYLJh2F8jt2ieY96Bh+ttK1n5KZJRvy9Cl1RlH8qv8pw6MRYtas3KZmYoaZGy1/w4lxDYyb1M
8j/d1txjabExDlU1aaBWaWeQBem6JRgLendNI9/A81oHKMS5sAgYdZCmLs2th/4tKY9KE0tFPLAN
oDBFAUGDPImHSxV1bZimo56Fw67Fm64o3D/WFZtm1Tz1phxm+X2Z/DEQUA5iFgeWk+2PZLELDHGo
7zYNJDT3wnodSka0FLLr6ggPdaOtRd9b0LuoPdETZt3J5pd7O9jrUp27YdTC8xzaoK30xHWaYiTs
20yQxpwX3WzIiu1ni9/iJLB/TQ1szCH3gWzeHRfu72UfnPnmSWD8XnujRe9QvhNwBC06hUcfGG74
aXpkGqCVsWHxbhs9tVGDdutQqOhjaSIPC80C+WlPRmeJ1yRhRVWrBEsxtLtZ0ikMWGgmQOBI98DV
Y7SEqQzn505KDkjIig7YdUd4WFJH2QACrnepLW1Mfz4mQhn7zg2gIR3bcxCewT3o6Yoabupaw7rK
+S1BeHq+APXex1SxApBKT4jlfsS6n9x8N2yvnQdp0jTJvymaRUZzos+NEZH+hsq24OZAkVJg1EDA
eT2CAmuLZHiNZ98RObLG6+68u3On54HMcFAE5fyNvqZAOO+VFHkXqlcVVP+C2x2IQflJmhLvcROk
6lmLDwdxDBdbgy+nV7VcDl3cAWDFj83ub5z9xGxIFsbXmhZXDEtPWmI6PSccCuZ+iyo5vCcM7bAe
CPkpIfMAZl9Jfe5N8ODHG6dBrhniHGOLZnNams7YItlUv6PPyhVZFE+CpG7htUA9UXQLsK/hh4k/
6OnPkeOY+GIn4iYT7sm5+ie4dCM1r6hZDDn/XoUR5CqCn1yY5SoGTf+nYWrD9cv1D0FI0BQ3tiM0
5XfRQqF2DesXRkxmC9tL65G8xHqi1TYCmW9Jhc/k+R5zdNbOVpIdg/oV6gPXEsPWuH5zO8B4e+dR
ozi+gG5mA2ZGDh9y+S5d+E1Rfa0An2bvPT171pJY15vS+s5nKjc5Ug+XMZREwJskScYkZ0EMInTz
J7HkXFn7qvFTI03EySJNeD4U49OfIhoASAWdesSwRnecYee8uf3mJtGyOToIPXhvN2eVGjfyAy1j
wCRM4W7O4oQGUNiGh8rEHRHnVlfrbKoMHNjncTPPdn8S8JuyH8MoDbPSagCn6adq+ltTZBcbfGqi
JEWTeqP5yXxQG7C9VXng1ERvbuFsYKQ8HYE2l/WRc7/5l3sRAVIP/jRt+Wcpov7rrDhQVFu8Sqgt
oKgp8YEZYUIs8VlTSJRT79WLTYjLbYZf4c3Wr/w54i2f9eCFvTxLt4qW2uB3hx6yQjyF7rB30xij
46hPMqEsOdh6CQ2ggfhDw+RBnO+lK8mNzX3tKKnkP0Wu147sglwzkZEskAfexbcuNodWq0cLsCQU
JLnw08coYQHYl+yIX6PqoQgNtimI+oWpr20ILYlJx9nMshJQ4oNdhWMHZdAPIExJhkTbHP772ZM2
NUrRijGKTVhYP8OdoNAio1aHavqfuYOSSeMnHk+jHp3ptgd9oz8Yzga+71yejG7edxBZrRDycT2L
HicbTYg+2pT7Y3woUc3M/m5hiYnPCaZh4au+VNEjQqSIJrtGWBrldA/e6jMDW/sSg0wIkBg+DISw
b7SjatYJNMZMJwNAgnntg2Iu6In68HWjgq3ebDMXTxnBbbq9IyN3lN/Ogaph2RyQruU7DZElPUao
FQlbP/6y1dFQG/wr0JQCJ08tGDaNRmjrXcqYO9qDD7NMR5+cVy5cQfsjMETvbGQI29ItQ5pcA7UQ
xA0yicOw5u/bTm05p0Ml23O296eR41w26B/Ins/FvZ3B9TB7m8PhR9WOPdx+5xJ2PEco3tU8boJe
W9BOQ5rXggTQWonE+GO3qTX6PwO4hGMR8GTPFEYWRaKAPdrMVK6YTbIRgznvPdfCWWvsj4cCmIHF
/vYyiJAvR6sxS7hNGnJIlsVDIDpoLtG+ejV+mYSN/oMxlg62LdpYVXfEPRMAxd7B9PdF3v0Td8jt
3BEgVSfJ9Utj2NyuAn5MvCmmJThanFnlzk46QOcMRCjaSvtXJN/C7RFQSHCuRyjv4oGf/CwiQkmw
pi6ykqbY0CJGso7RNsrkGyn8mI0LVRCmYApFzQxwcgaGbcPeHDPr94GZwiF8XU1bmc+S0BCTJNkP
r20aNXScECYnUOtJuHhRndwPw12SYJ8j/jAtoF7UyT8dyC6hYHyOkwphsOBpkVXr/nfAPtUsiQ/h
sDj/doqqNeqybTMEch8jdICjf+iN6EnN881j3KlNozVJ6XGf8uLOi+uKISf7Om33nisFA+DeTinP
tw3kJkW4xPkXYJD5SwCBXOJlpgS1wuHQMSrbkzE65zFPUWQkoLH2u37L/dk4ktL4uuA8siutxEAn
SUUE+Gq4TKjnCYRqlQ8YOXC82Ni5lWB6HGz4ZBzYkDB0FoXn5bxybWNRSdXyjZhpLXGYV9eGwrBC
Q4b6ubBWcMwLwHlLSLW4szFSdiWN8pg84KUeVau7VwEwhkMu9kTsh9BXT0jNKLCCmMbK+Cy6NAd6
0mH6lmxqPPykLwcJChRBnnGhti/I+G8V3GJiIDGAkNtIwKljNp9m8K96bmdBsU/zgUmM/POe9gBY
io2Ida+GIr1TanAAET8YUKsDVOHBqx2DZdxVwNUl4PvZouDkgR9TyJFQdiDQB8q8Btvdn96iLEpo
WCjcs0ShzNVm61rCHQkOJ7DLnAYW+C/JYrz+CU44bI6IsKpg9pQgQYnKynnH8XDpAgrTnz401x3S
0gsePthRoUpfezI0NFuaqVK8sO8mdE+oWT3sOjlP+FBsIFX2800IWXTH1h5wq81C+45AJyostSLr
qCpjESSjRyFs9HvBAQNvIHV76SUrFpZZ31PyzCEDRVl1LB+DbEgw+cFhaissFTimGxuQfWUQpEh0
FeF299GOvYojPvPXLo1vhmJhVHBU1R9NXYQKQT1qegzfYBb2uXKE6i1HtTv5UpRx6cxHYCRJAfn3
oB2aMSrXKPFh9jSl6KVZatJkYwIg0pd87FbN386oxbJmxx6LLb2oWt8ucPFrPa+bVEEre6DQgsWP
FlHz43V1Jgs8IPL3pQsNGUk8h/w6g1J/bUX83Uvj1m/raRgJWy1ba6OrYHx0U9oZR2ZXWK4CEkCr
/NA/EGEk2SKKLG0v2vOTH3XvTfrlCWJ62hY0/077ZJxSNBZpwI1i7Qp1rVkpyIVOjd16Hta7O2aP
suILW0iNHdpPxRA90pmCro1G19RU/Piteh24GAbjkC8NUbumhYJFKKEQKatqtJP7HeQVp/DBAMUc
mkqdZbF+QppvftcHckLO+XF/HRDbnUyZyRNeKhQEsbYtNkt9vs7GCqy13kealLgyEJvTWganM46M
uZqV/tBU34Kw4FLg+7hxbKkpHIrNRTWoVAAhxxPxVTsjV3QvarHCKcBd4Xj2XQYyWmjyGenHYTeq
WNSyFBQxaqO8IZZHDdYYjUQCJU01U/PPdxHMUOrRjD5It9BjqNn0bBP1/6QZBTRpHZNAnwVk1LfI
Kz/aKIQ6pw6Ty9ebLoaAmtkELYUiO7QGTJOwLwaFbZcoIH5P0BA2lqqBjC1o42gGGaBz4//6ablN
KsivzS2j5uxyFKzC9nkGHSfUUoLiVK4C9j2e9S9FYb6cB+MYi6X/WudJsIeMYb9hSXdDBgWIOynZ
9d39cLRptPunIzdfs3fDJOo5fvvosVfTTZQ2pbwxr4oYw2tpGP9NAW4Ej31V/amJ9VARYcErM2gd
GPiwscFaKBMt4wvnouQ3a2ceOQ9BYgcXLuq01+iyoVoYnwRSdeU68cYtuyjhvCIAzkHF+vUlv6rO
jeELSUHH6CNEgfqDL8GeTwqd3LOPj2X9g9CKrscr0U2rQlVqAoPMqbuKqDfHu1IMuLqn2Sd6ryHp
/gYJBjJZebyI+gFetgvhA1jgNLwJEgclsPAwqa3Juhxl5mx8g0fVSSciEf/k0BpDdgZWEZwbka4y
yFM/BLiHRSQYQYcVTqA2kbTevVT1z5kwg/Lih26kUZuK3ZG1CcelYn9C2T/x7yG6caW0ApczlirD
eLxMZgdslJTP2EMhQdSp+HNkHmlirndb2F43p4fIa1v0+FLEu5YK5hxV9iThcUxCJe+VVyvQU0Ng
d+RkuFOwBQOklsvKsp6ubpIORVme/ErnM6cpmu2v7CdhUiY8QycNxJSCarO84jhUNt7ziN+ltaKo
BWVmzKRuGoXpBBnSqxdUCxDeQb9XimsKLhmtCGKul62d7DBvGEPJFZfBOGi0k7zKlX74MWY268AJ
Hvkbvv6UpQsmIzefo7O0LTa+sP7r8oRewIAQuSUJm2TL05WDCvDYUUNYlczS9ot6hNsfZISfZkIB
ioAvq6wnKfbI+STjQXXsY8UJkSYPusjSilIclsZ6hMo7tBPjcnfrhZ34WqQdLwSEQys3ioBVNCBW
sWNDZTy+y1hmJ95MpmY8t0Lk1CuUDI5hwZmnIN4f3H93FeRHY1cevtOtzyKVEW7vCNRj4sXz09BH
oWYL29akSldcOpraiLN5vuPXT1n39VCONjFtN5kTXkMY41yXtu49SJOB925+Ly2MFKcZMU4F+Iak
a7UKhu+U+UjJYprQ8GAchjodxseUSe2wJ6J4kHce3shn2L7KzdKeT9S2CsEqW5f8/GyEPl1sW5yk
cb9YfBlKPn0Al8gpLOnplLDnMj/B1oTsT13TDbvAE6yVsU/dYYhf8H0q5R7/n/yHjOa4IwtaA9fc
9hSFd4qx301iBOzdRGGAqq/2F9+pLRaBGG6/Spq9POMFzPhjqQL+tv6uhva5AEksYsqbYFiQuLLy
X3V8p3IU8TWf6by/ocL41fA7C9thzoIGf936QPog+8ckv1eqyZy439eXh7U+KlEp8/kIawqnYe3O
txfjFQJU7ODDcau3aRCtOwPHIObPapsnyWlpeIXMsaU1vF6Pv6mw4c9GPZSx/vxRVZcy8yviZ5iY
AG1c23YAH1ZJrZJ++hDIW4YnOHFr+6E+WUoZbin5HH0nbr0zqQhLp0YllrK2eJ0h5lriC64k19UB
mQT3Cu+gVEt+pmikQU3UwVt7nYrz/TW9ml0WISHFou/UxNrjNA9EqX13SqRpkRknJrfY7+e+gmCk
eerSNgixg69T4s5xEW4Hzk5QH3vmoeoveG62Fydd4J9g0Un2WoQu641y3BYPAJ1qPFf5N4AmRwSm
MZexfe8MEt5VSQMAPzX4qhBlEBv7bzkErsF4pk+nIUYs3I1XsC6ALwCOnAgdgOw9jB+32mZeKUTQ
9DOkKzt/FymV8NGyC/uucIj3o3MPgY8s/oabgMYo3CHOa8hNWZs348cOQI1KU0KwixSXst/E0A3U
HqX8QFo0hEBB07a5jklEXfxpwxYwEumyOQZjQq8rXLZMUPuHJNmc1nsS6MPyfykbgWhSJ1xpfvTx
C/619AZVXZyTzGhEq8Yp/FG2+IEdVaeP4OKFQdjoNSOpn9kx46HTRqtq8+i3css65yphd1z4KQNH
MnHjrznJn/ejFU0ZvRwCCZGg/ItJFC45zg9ZE1+MEeRnOHyOvSQpHVcyizz7Tc4KeZfNFzKAR556
XrdxWMydomEw4ZQWZNnKJ1bN7FhQY+X/8mnaDvtFiqIFAEFZJmaodTYMkneiOH5sMAVL5JiYMWSs
+h8JzjYRRpqLGHOgp5paDgBDJSIh2ARv/rZaRXj6wlhUkKL+FhE3qYPB4p++xN+yapVfQWfKagte
UdtN2Ipcx0FYIz9o+JntOb44jGCx5FoEJvaLY16hrzzyCUHNeOxpipJ9S+17EOPAwyrHSCOQk552
JnDu8d/+NcgVaj5bolz7r/bEggPqUN7LELbGNy7ATAT9JqZs+zAQWF1BNCt1Br5UHCQ1bCxEH47P
vkDLVr4nOOStdCC6CWBl5kc/y9IBrMKhXoGD/XIB8oBN58OaWmjyioiF0QLIT6ju0KkTLg0lkcKb
6QSAT0+uKliY8gKO8FK9Aj1gEW9xWaWe59nm/elWpV6qHMXJIuqNUUkYACD0Z2eQAL0KpfFW1Bd0
HPpNaXD9chr3Ni0eMvXnRQEmW1eX46rhJfDHya57yrSFrVigUkDN0J/q8xPjpbdM6OcXpxgex7+s
bxR+iIOnTV32PeK9StjkO8Sc0MSpYjPmJPgtOniGvO7SxYvVv3myT6FXj0FHlUCJHx3hKyn6Z3ae
gJ1F42YOcOlBpwhn3QYm09//H8CmhhmG1vLoiegQt5c4KSbS4dkJGyZJr/lBHiKGmEXPeJxYHwDf
LMRNAcwWvTDO4CD7OkQEZEG/LRzQgwH163B+xQ/cJFEKqYpd/Tb5H3cUMtkmmddI6qVY67aFBVnh
t4ALzMBs2QkvIjRKJQmLUWk8u5tjP5bjV+/5juTv5Rn3mSIIx3NHQEyQLrMBoQfVRZNmK5YXhuG8
ELRWSq0n3H2gyJybunorqDVhBEfGOzqGf+nawBsSvoT6/YfR43L4fG179OVlgPtBZ073aGMk06vk
53N06HjMXCrsOQE9wbpe24j4KcHgu/ssYtVyCTqhulykKNXUAJWteVSMy6oaRtR9sVxc8K1BnWfB
U3pcha2vDMDTBbtKU+xWC7/Q1osWbMdnLGk9LkF4YGZdRYrb14s6E14EVYV56hY0LuF6cVLG4F8W
OIQx1rTB4g+d6uHKfkYnm36snYpOCUztIK8RCBFkPuffOCoY3eoPaV9f3Q+HkeQsn+5ANqrALdS5
5fIAGIN6ziq1czQTluPFbEVX1OGpYpmHrJ3KrXx7GmPhQ5DYO7GR/0TZhqXgNm/Hyhduxyi+pvbr
RXVbDN55Toj2zJLNCCkPBWKoIFrBiCERoT86RXS93srRM26ZeoULStmHHNJuqpVFyPRJDb4D8OmZ
L3UxM/vTrwZ6g4A7CyL4xrpEJ5bUI5UdJjiGxRc/xVpcnbQMjNtwiRRgYqTY7vMmEm/UPwponA/R
XPmNJkAxqHz4gWsUqG9p7oG/ebcg67ZJDeGLRU/wZFij5xr44hOeynntdIFzYrRPWr5mXRycNK4H
RsdTAu0G5BOfwe38/rba7r+o7aweWIZAFsQ9jWL9Ed/cgi7V/flz9ZXqIT25LK9WJh0RfztYioHM
v9y/CkQYm/Yy0V1+F+hSDOqeaTp05YfJbENsOOnCsiqKifQubOqOK8w5m9Xfpp+HHlCa6v0o3XuL
3Vx9QYUukDhZVk+L3a5/Q0nnfH0xxrkiuLgZzsBvJ6gwfOukiWtVA4gKFOlEUSyJrjxM36Jlq8ti
+gmx1pC4gOsI/6X9WUDEkKQb4VPoAu+fTesAbfce2y1F4dv93V8CO6PdyZBFvBsmUVVNRkHauCsW
fwyIK2apm0FwDy7AWNBscHmm2qS3jx6E74I/0lIbRTLVAB0lHHPzKt7dzaO9RqeggydaY6rNSiQH
OOG99a5xqxiOHHwjlbR60JTrFc9HVsuly9yuH+RIp8szlnkPaM2y/Jv5gvdexj3+7o8YRfFLhSo/
rL3iqAIX3jbrxUbKGAbQ/x+NQoq2df6lwOZ7x4Z7c/g0ayp8hJ6YKzilQ1rsOxXqXZ1lSDFYcT62
XGXhv8fMhSVMwdQwcSqV4pTl17+XP2K/IiQhp8oxKxq0QTQ7jQVTsVwchlwGPQS3mZO06DtFSl+L
LR7Ag3WvtSUbUiJCGF3iSgjUSJHC7itiE7Ap5ncSwr5ontXqbtFLkylloAH/JxYLQ54Yfn9Iz3QC
6bnBv1zk86/lnCfKVUPi1CVjOHGF3uIYn+ZFrwKE5cJujNAWWR6vBXY5Mhuiq/d40kaRkfWoLw4z
lBTBn1sU7WRqXVoNhVrL1flg/GOaLweMF0D8zVWVKQBbs6v48UAIy2g/N05/Bky+TU3VyZjfypz/
uW/skugjVd1r84RKe1c2LehTfy2duJaUCgOuJYODrj6zz81lCPWqi+C4nAtv+ua8qoViWpcZQh0z
N65JlfACbpNOHwu/WvoNCR1PrLamUwHkyJzYkYKDJjmIEC5MHsC6UhjZhqkmlyMky4wg+lG4tZyV
I7AoHEv7G3hjBZzcXmY7kZ8Idc7t2yTP/z36QUr8THtXALWXJhmZSsXswJcyzUCa86gQ4xbSz1l/
nUibDdUIKMm7zg4YQrujkzlWaFG1AVQc0hXWpdRvwTYV66fFn+7las9eBw0cPRSUzr1ny0qwnUke
XGeUVP8iXY4Fb7l5PUMpsjJ7Po+vDFDkmi6QKzURG/sYfzlJibhPabm0axIOgmtWjJkeaiZdC1+q
lRxvuyDqhh0DsyeTkVRAz12dHR/D/RHWIqzvmZenic/KX1RC3UAuc76HT4pqleT0IKQLOwK0YcAe
oaTeH+0L3OCOY2PDhzF4mrBl9yX1F5vmyJI71dGA4ySErG7s6Li4Ab0L/K7T2Hbr82k814fPS1wm
Xxa8VshOuns4YnEwXULuFFyxiWP8SYLmBiqMvMa8uAde6lm1jb3FUK/yYcufBjQCCvLs5FysA4k1
7GDFLbr0pYIVqxRVRIujrYKdSll0ooSGG4+PGiBqZBqrjygKFlzgvxG6Eb+uV21nmP0A5kJJRiHS
6smKvz9fRNvwX3nE0cSF+b0qcKi9bq8SP5kLliW7jhQ4vmbRzv11rfSd1cYFM3hIgk+W/wTNwIvy
RGE93qjfGu82BsnTRxJNFLVU6welO5STtaeUjNYXKd0+X5g6IA3BYDBZWVPiN6Z3DT6IPXXAcCd+
XZoL4KqSCbvLtnUAftQsU6krPMYnfZgxXG0iiA8dHskh3mUbTSzFcPAGWm3wd4vn5YuE4ONsIYzf
RyI1DI6brrOijJTBV63DIPZb1GsjoxdwSVw9qlzBh2MAmWmyYOPhjyNIgy1vRjaEXa2SO2iDgJhf
A7SXZdRcQ4XsalS5mLq+Owu0cyWasnTlRObYRpeqxyftcDYxQ42XQ68i+6tv8MGXZ5MgdazjsP5e
XB8nO78K/kGFPhLaoJ/LW2ZAztVz8eKMPuwKKiWMjHJLtOjBeSLAE9dJDDbBV2bxABecvGAUfm3j
JrZCyTYzAnhMKcwi0xR/KbgWqrwn/fiRNbygqXX/wUQLbZQOm7PWUIvCNyJtUkmXmx1jTxU9a2GO
JnLmIM2C7Tl3OXythUWWEv4lONGmkIjunbKJq+X/8OwYFdvReN3AtbZKUiVXNiB0je/ghJ6v67wB
XLyZPmgqNLQ+NKsoiwY3u0754o/opzTigQz0FFxah21oQCdyO3d0jYiVZXu89H1YFOMDL/BdS1CW
oDseesqzHX85In6g6F7Xn6gnbGYivAZaaZBvvIj6HNZQ1S4yU4/VoDhOBnUfs9Rn6ar2g8hiW5GZ
6ql0dy1MUSBZg7FaOqizVQwIzmkmn4f+pOxIxl3yA6DOkThjg2110GX92lVyuN+2e9azeCPRezrc
1S8bnJThDG72qZ1IV0jEYGSQeNa4QmlK0Xy3qTLNkHm3z3fHHUOkawc7nmJUCJHWjwX/V2TZMWF1
pdHs+Z9/OKovEbXjxMzobmeoNoemOWkA1A8wSElxjqxZI0jUdEaufT8F/ErE/+aV94Z9kloEWXuE
K9j4RCBOpRN3/L3wyNGTsx7Yq4KW6ZJCzTgF/75Qeup0ky7ku7m2E1QyDmdtgWDiwr+N+1WnftVO
WUKfLshoKLLjFHIxPeM1v5kZU6AfJ6VvTA8+pqnh0s+WmS6IjKgb86GoAloa2QtS2NgWnF9xM0yQ
k+2qZyKfn91eq2hzKcPtmmpzTynK4WV05/yNOhAa7mMhTWfiDT4BVK37jRimZzf15511UykZwif+
IghalDQsfO5XYTxjWpV2VAb13fNDII+4xIuTgSEiyfIubUIsRhKnVzxvqOAwPw6FQ3Z5yCasFiK3
nhKbLa9BEJw9AAwEvTK3I5csgvC88s4ZNDRfPXtipHoLsDhwnnqjdbPbcZq729iTI89rEoNZ4Iic
trjB0RyggGEEGVca5vAEHnN2eLKs69CWwHkP71oTt6qLvjBdO4QPgYyAWwoNwZQMLqsE1IXwmK/u
YfVqtAV5wHcJUua0EUy+im2NJ47yzBdtcXV0t7x3QkF7ROsjLkiYKp+heLp2B0SGeNOUf06oqTTn
A/FeMP9UsX9sTJMxM5IJKPiMpvHFrsT+nnW+qGxbWwWK61WT8vHUFRVLgsea5gP0SC8D4n4G1N4T
Qze2NE5W+aPTwZYwezgtSGCj1gqmP1RiFqRBGoRwT9cdIHRlg/ASt+ClLRK4knOICy6YqpvvESWS
hbauv6UDy6x15QzaR+lk1KvW0kkwe792RnjFRA1l4utGny66C3X8PPtFtoN0HGOFDTkLb92nnmut
K+/mzp3jPNrAAm6w7UP545UjBGvQAuWhQUBjP2VhxgGwTrTJxGVhOtCHiN439rbjT19eUzzy+zY5
2KDCNxfnDpsjH+ILw6WioAJXVxft/4CS1aN9H4Ox0jNVabrbJg/3KPu/SdbH+a9KUe6xbixyfCW3
9zfL4Iv3TtkVPq1s313rdrbAc4jTJ3zTta73gdRJdnTmx+sOIrtintDeXyJHB9rNe7WAOvGm6mgy
48boIWIGyMzyzAURgI0FDgm3UBLltwIIH1h/blsZdXXpZTFdvsyW1snHc5fZNxWqRV+DNsIM/YJK
hVP/iKUZGRbdjxUdK/KtVrB9mPQeExdC+OwW/+LjxN01++CnEZ8x2R8msBH3YJMM/1DeYKc0eQ1/
Oc6OcWJjXYszt7lMaTgwnbrVivpWYlO1iorvuMA/z78zKg8BJ2nLP3m4ebdsKcd8B8abEGZtqEVt
GRFZce1rTWqSra67bRvc+IALBegmqzQcuGec6clRQLA0ha8k4IDK60wUMsJdsRRHPaWFja2Relji
RrD66g15Q9BmP8m0fsr8p50BPgVHno8mKy+uwHuC9aHfAxyO5Zkr7RXhQhCEFBbYrBL9th4lvUwi
SkmBbhms8yuL+OIMBZkvatmc4SNRrlL1rde5LcybHRNEJ046rWZoO8yzvGhDsWkAenbPCaOfQwFB
0ab0d5FwwzaQcooHl4jjdC/HftA6WGGGugiltVHxMK2B45k2HXVR6KpHw2ZtrUihAT/d+7qH/Ta4
ckOmPutp5v9PWQneJp9qu/YQrOkbifgmtGy678CJjUNFw+zy5MGCbl171d9B0v82caERlvjJfGak
aPvHfU6kBhACpU2eArwCxq3KgxGE4wSrL09sa1dTQHcjBFrPOT/mC6e0QB/4aDdS+v7+QuqHXr9o
y9hLF+Mdo65+k6dxTMNExF0hlpVN9FQ6jIeR/C9KVvU9P5iea6YCl1rSgCIgVBF+rM440hJMqed+
BjbLF7lYi/FJ3OhcXDbRXeaHuXUQ7eynW2w9gqYhGfADMZbw9Z6Abg2ntLb1wHuuS6zW+69gnmNI
w7ilqn9+qTes2btpd8/WgquVdwutdlrjkRT5sg+j77g66K5V70bIJQn+kpqlPqq0JfRKKHEeJbcx
7VxNMH4GfMUJTKDjgddNypLyYgZT05/2eTlju9DEcRRhAgAFiykFMgVM1CH2dJlVRfVeGPWKsmRE
P3XHnqTx26Q+TJV5Km+ue/n6HSDWFtmVAUOAkPAErEwnjmQnXMQs7NrkMBUO0ZZaynS/QIkzW4vU
1ay8UIqoMW3YFeimhCZOnNkg8+/ipnV3apAi2h7sOFfhnCDrv9y7MeWM3OvOR6vgqN7nWJdy5zTG
djaOhg40pVbL4S2q8SbxRMIKFYs5q2Eb+yhiRF5LTAzfko5aebAukCAnMhAEwEED8qE6cVYRj4jV
koktfuTCdA2xhCZigG0u7WJwSwdE5USRgcKW1iVVxQ7V7VfmtxScBLFFPteJdNaYLD2WG6QV+gEv
xe0Olc2PNZZVY/xQgSlBM6IdSz+4c+7zrcVorzdgKlKJ4Pi4ivI5W9mtVCtz6Q7up4QIU22zP/4h
iCvsicKzGKpZwOqAFpmWCvSbDcsFtcNfqhZ+SllyLD9RVZY1qEvs79E0CBp+7Au0TQxHRBuyrWF5
58JE+QPoCupRbYp8CKxuuLV/JDrotMI1aiIcozpe/8d1ZoThrUIbjLHPxOl8sOCYIDDnhJ+7jvfL
6l3hzxH/qft0OWYOHsNRf7sEtAx0sHUAjzVgtJ0CqWWT+rZ70CLLyILQVyawCpnjg/Fcp0vfpfmo
sXD8ChYtfRA5X9B6Mv5XBd3vKveNjYW6XjfPxuAEMRoOnyhYT3mukn8zi+YKDuWhXrJzEhk2LhEA
TfvLSG7LbOHEXOP4Dj41WpsfPvifRcnLBTgqElKoHTJ7+vpMdjWExcADQH9gs0rY93XxSsK1tIG+
0Grzblr5gR6SX83iFKjmLbDxRetJg9YNsXDSP/4WSaVTuyKPnmhT872hjWODLf4Np+eisya6uMsh
aLh77uBlQpoRCR0bjQfYg2fQONRfSDqEjCTIHSEN/KwUhLxLla+r/Dmds8Q6cHURTqu5n/Sao2cm
YYjxXEIQRdmfMjTDgsj+q6WLZa/mBMW8WB4+ZsUl8XyVrPKe7PldPeHxcLTav32jhY2tVlHv+hpk
5KfMj+3XSk7Wz97LQ2SwVIlMcWbmOrhLbQfUqCy4f0xhYJ6EB09wqhgV891UnuA6ezGG5NRVrEKq
5F6TlozSYtHyPn+lcBYpNNdP8g+GxxYFrF3v2dJTQhf5ScdZULrsyHtPvhZCpKPx6tOvjgToAaOn
Ja5/x1ngDjCiQ2mr6YWRMUghRmsaycyDmKwNLJDv8btL34zxDUbnfAMRgbSwj5idJbmzoOOtrwWq
HWrfaZfaPZokFBQPYXM6yH+tM6boIMrBx4JIXrKyY/xI2mqYFIWgLvqv4HaSJOvt57Zf+UVmC+Hc
b//Rt5aYJhws6Cok+xrJRcIwLLskuZjk4K4Ym1QT27c55YlqKQEdwg0zskJSy1DGOzzDQ6SHSHgy
u5sxEMkBbINpqTRdQIo7sjkXeXRh0aUQZdoW7enfaPCwy0QCrtPuOtKBUP7lH67zj3nGvdK+JTLQ
Sh9BnSP28QDhY9tlqBJff4yXQ6djDSj6WFSlLwH+PBAqGeVlzE/IPpHZP7I26lhY0K9DPSwem/W9
vG5HhDlgHrOfcJbLyvNuvIR/GfoATdW/9cTjdAD1olBt/1YACM2sNQtPSI6FRrXbymveYrn5+nuF
bLq85lTamM5IVNdnEtSPARhQQuua+Or3ChJPSH6WE6T+sr/RZ/gqLBQ/SNtD/9LXUV9j/qgjWlkn
IDATNawwe6wqU+9LyPg5FmWOipK+TRIVHlkXBftdYRL5o5KtUbacnDbnCnsh1eYts8+DuNrPnzyd
8bOdaaiJPpmyFDDd0FFgkMxWwpq7/blIWKirmxe6n8shRoPF21FGc46MYGEYICV6me70GGCiep1L
8NdfDTMM0Djz+Ef3aSzSrLgzcdPlFwx8YlOrxK7943JrFwUNGRjIwPoaozbwCqtCGmrlCX0bz07d
EX4xb2OI02AU7LYqAmiylnJjQT62pyP651ElsBH9dptEe1FwsxNhoS7NPP91qLVePrGM8Pn5rTvw
xWXswIOZh4oksUl5xX4l/juZi14bcauWprjoNtxNXlELcvk/GOafYyRBhJKhpX5P9PBHkHFvvmjj
wPdk5ePZKWGXump3PDG1WlnhGxzm2Z98zewY2IoZ4FtTYHOuj0omaCyvffEb252sBS2r9JadQuP5
fPsMXc5gdyGwoWLJiy1drDflXBgRWNUmYc2cX//Ted/UowIpFsDSwUP6711Lo6jXHR7nbx9V8Unx
2h+bzzhpuu8nXIHBLQdrJhcLZ9im5f80aKOMPJwQ3E1ZdH5JRWS2oDamHAYR3ICbmX53dAIIW+a2
0HTwN6QHYdOi8M4ZjhvJw7omcwt58J5wCV3ai/vGWN4AU//T3TJYiiO56NTCjlVNq+wOe2R9wWwv
PmcqHrx87uk8tH7yfw/YD76uUIULRYa3MHBXVDbdkXfvDnSH2lJwfuftyr3bzmEmgNVxsL+3aQmd
QKEwbIfspQhdC9tCoJ7KeiwyxM8sT5SYW8k1iU2ymPQrEyPIGfOUlqvyoOE0tDlieZON9q6y3rBc
BlRFO99YCdtYU1Db5z8iiOlCro4NTHrm+9XWk+4MtZm5uyPuUbwwRoq877iZ957/rtZphqqrzuMY
C6uM6H6g40ok/mXbVhy62MK6tONqqLgtcIUDISMhTkZHQjBcDdBxSyTmMcwOeNkOIvvKXyrITQHK
owKSB7Uctll6/Na2zy3iR3WmK5gP/6wyPRxbzMz6iUg2x4upCa8i16siJypoBvZJCqeUQRnh7kp+
M/nB9eB4FecV7QTMOdtrALFPkW4hdX7Ap98O3r2F45mCSYG+L2O1dCFlYc5Y72z9PGYnogkST9nm
zDB6ac/BrSeKkcHQdTxHh3gqghicPqxQyjWRF+JXr+KJxz4YVHFNCADZjmvHQ5pkVnjUD0LR9CQM
iKpeJsuj3os0D0iKJYb2bDbjYXf2oVovdkZfsJYJoVK6rb2Z41A2IxmjbrPQ8BKufJfhQPj3OlyH
rIj6brsH5YPhTL8B+JzpPtRlF5ALAKvVcnOd94RLq+p8y9zPeXWgPlcfvjqIAwZ1NM4awk2WsM+y
Py6fcceCgz72D7clWgZIamNxiFb+J4CfYI6se/Jvd0EiZtZfUCkKvSdR9evLxLfY81r1AENYea3L
dlC5NWrmu2oqRJObzeWO2KgU5ORac2i6cMjXK1Tcl+AVbhfHPmhZbZg7J+8WTEzfaWphKsu0D9wo
QUip43sSNmvFrmENjUZ8npvU2uav71uqhtoskxCH/9ddblN5bUPoXOgARuBN/FeaW1eEJyxhlqQW
eaTc9NBv7zsT12rskSgmCEzG4966pDR6Vbe1AyDtgXuvMunX4nmJljKF1XpPL83wiRQbAWJjMSHv
fxW8M7fe7JMRJ4g4XjLlCFVUDT9clrcj0W+KUVids0pK//xFpxroakAjqguu51fszy6BDEAP2lfo
OZtSGJ4yzXo9BIvHfe1wtXZxpBn0VX9/T7AgSDA5dIexwbYitfQfM6T/otBF80SA2b8v5BypwLZ2
JbnzCqAbzgwokAjkDnk3gb46au8C9fqVOX2bSt1yQOjFe3MRnXBVeutdefhj91+Zg4pxVPayCtwM
pDDa2btW2Dugc2H+Ccx2VjOMCxOfA87jQ+xLOOm3gyWLP31JtVxk5S6eIoGa7FCxQBhsNBY6tGet
Crk62EdnyuDCmF6L48LpLT+9CO6G3NMZIClXu5eiyspR3XM0u9cQpS5xvDaI/JX0Uin1KO7bxmxv
gp5i6EfWnE5d7ykm7CFslifsgkO0L6CWJrbVgxiSabenptAs517oZMbFbrpbB9qA7Nf79peF1RVl
l/Lxr5rgsWGpojf+/O4++2VT0YlRZG9F3diR9CHp0sxpkbaZxJPaYhyhD/iRDLkJIHUxgyYljrdd
XT7RBK5QbrOSZ7Q+WddeqfaXJm78WLniXAIRZTHvDbrIEHZG3aIpHuwxoRjraRXWDf/Kpk6mogPR
m0LK9w6PoTiEcMcUwfHeaWB+2HuRuZZo8H4s8Cmao9a22Av7c+fpcMu+jOSqbOuOikUEcbu4qnF5
Mg45oL//0qBd+ci7cYeC2WFH+g+fhXL5F3IvbAfM2BlE8WpSQ+BSIqTPxxI24FZ3tJBhjkZBABKY
mgYXj4aJwq55SkiSyFK8dOIjJkDxZbEaLIdLlt8+q/p6dGJv/b/UG0DVkEI5gdrrMY/WaNY5mVjf
S6zs9oObhgIZYldcRFwOlqus90omVI+Gc1dDdG8p3NtHV+3v9ZJV4DQYzkzU6K2nuu+hefuxRpoP
883xk7JfDgNJQkGXfMIjEIPERi80Rc1Ml+Bfa5e2iPbdRGXk3yfxSeVGc4NtXwHNFuNgccRfhXBh
SAZWkjm80soKAhzWhLM6+8MStuFVZs6t3m7fnvM3dQ0P8EyKfZWMJS6ro09w6X5QYkYL7Yz4ZsB8
c+Yee0DNng5Q+KUO7h1lKzNO5UZiscask5zZ1vir0wQf9pwPWxkbT8UV7zaOQZA4QB3w/1BXpx4i
KuG+o/z9ix8D4HJwjWTTHM2Ccy1/f2v0um3KZwa/AjoZFWj4P8FaTG05YzaEtJ6vOnXc1OTBOfMB
RyTAXZkWKciL6frpKrMElIGWy1MgiyjXPpzn6HFSJqDKS/P1KtqS5dXTCmXg1WjoOxzCQFyDXiuZ
cVedP9EnpN1hvYhytRhiZp83StAU0UVgubdLozQ66Cc2CC4OaH1r/H0l2dB0g/WQ8HzpAW+gHC48
9YaPgKV2bGGkpRNK9MB0HI94YraBFQfYsGa4cFnxVsMCILguh99irpj14pJUlJg3AT2fLFGRtg2m
/mHdyIRaDGUE6PzzMeaAwZBQSMwYMIL5uqgtlNFIjuSSCn6lKRwo2SxCZlVHgnAZOV9Y7SWDANFZ
lAcEc0bGANrTZPT09WlOb64qS7qQdDtH07S5BjUuGA0miOmr9sN2IP2W+wUbDe8mpg3mLRUWaNT1
Cir84YFMlwNomt9d02FPdayB4pfyi3DaORI/oRgilZIKg3z+USiqXFoc5BHADTlwP1bVDZ83UWkW
yHYVOuE1B+LWuysI56lm9NBTvMwbBLEgm87I99CDT60TXo/Ywjlt0JLqEXZPX+vszu8F9Nccnwjn
c32GOD1jE9VLcs7vTOhS6bl+SF3dZeeT3N/OcTA0CgxmpbU9Lq0zR7Llk1vcT6cPiJ8wRtN4JKoG
zilsZqVO1ovm0ZqrKFJ5UR/g9uAtJgnId3IW3+6C+lAbynco12vzqHdlrkYJOjqmi9kQAU/xRdc9
3SH169U+uQJczU3CaoDdzKGhEIIuBC5dawwRK3M9m+844xC2yC1ftIIDJikvGkSp2iRcDMIGyeI7
UVi6LdYuZhMqGhtM9NKc6YCMKpYLBlQx9ON+f77SgF4ke47IZoD0sFycI8pQ+CrtYqIpLfSfPVDC
gTD9rDTxqMd5jcQbfDi1AS94bDBXIzE31PTXIzjycAQLEmM649Cs2YBiemsVYfSa/X2BUovnndkW
pEKCQsE0c4yKEdgg9I1jnpmkvf7E9dK0GvZRQatmkvyx99r09NSqaV7lniZNLb2Y7VSovRcmzI55
RSMDvmIPteNxjHUQBrIcOSP3u/l7d1Nt6/uNS5IWZ23s/r1sTpkLIUO+J1MU7r7pwZSH2+PSrrQb
RgMqaaWS+WfcY1TPpjguUPmjvi+5Hmft2f+LR4F7ulgFyXKEXFlAOkQIpMLtoXVF1+SsIyHLg7Ik
hk7ctwX6qTEOcs/dcL2MM6FoKX7dEi1iUtclUaXabf69GX26+u71yqoewVn+RJTddXCuhgxkd1+f
SUx7NSzbiF3eUO4v4GUs2bOm09G5I0NRU2ctlN2jMvJOYWje3SCYCnXa95Zo4YITIw8WFgcvaP0F
HxJjPBFuI4YiuYaSn72/P4Rv2rskR2/rJ355od7rFzX7qCbDI3F7gQ99Sx0YJ77I/ZXf+JmkkZuF
bq/OzPGxHxZXJ9sfzaHQpKuE96T0Zi6g3RgiLJGWug34do11VxikpbCFSLxeUJw22Yk/aC8IFGvi
G52xLNR6YkhH57dz+J6ZJftix6z5l/GVUHCgFcaPI/ryRM7oVayF/OU78abG30p8vsvIoSewDqMM
CT4Q7IZVksmjumsHgjj2ONQTsLa59yIclbwproEeyS8mtd904Ar8fFy7RdLjbKhH1OEn69uC/RcK
N4vxwBDU9XzSB8UULS63S3mRfY3WAGLxAfw87NCCu1zR1n5t0oKDXo/zxzmaAIDJzICmSHQ4PQfb
TIuHTH1FhPacuk9PPX4eoBy16Waykl0yusHabPutR1AI34hSug8/qPqYS3TLHXZhjejupYgZ5oyi
VI7pNXVApmVv+k2zD3rMUY26DnuR4GopaaP1KHViz+A9usHIMFhIj23m/oqhW69aiudlO5o+etZx
y4d0msjTlbPqtNznyBLb/2rnRhtfYxl3SdcKOqzYBu+z6TAjuALpkh0F3Z1ycRP6XTWbtbKYwrXW
OJI+pT+NGTOmVrCxoifa6G72hf/d0+vAyDHgNyMep8e09/BBfz6l+XvUpXw84wh4GZZadWMzr+gx
ZUzM9qnPt3IW5bEwNB2OdWuvd+tpx8z9ClYTDf/KkFzCO/LgaaSMEqAS08MYTEUv3ZOCoVgdx+ks
wwIevduqdqnlMe4/InlPU4Ueo2ijX4vvBLFAo9w1EycUxjZAeDPTGeNSXXZRP5T8idmQUH4bZyBT
oqj7k3zP2SOgAXaObRpPmN1q4B4DywZXOhRJi/u/wPDag9fqMb4bWLw+Wt0TZmvP8ivrtF1AAdxx
6Jk5S8JWQ3SngnE8FHO8sZ4hCeOiVS+FDkHVICtrGIDICwAn3pOLKhPjB9ekM1TD+rRKGwrWRuiA
K1yhIMkOmSPTDhkXGOUYtncS2Tpw96x1v9ne8qKpoEXxgWzbrKB3yIt1CQiQd4rve68hgXf/bD4g
xRsuMhKUsMq3CmjJsZMNahyiybxo4dJP0vxs4seyjODxS5OkUIsywtt6AmjaMIZg8dBp312OCr1m
5sRy+MwBDTt8kUZ+X7ZqeJWTHDqiCcLZgrAA4O4zDNvamtLJ/ovLY1W5oyFG/zVPd6l9GuMOj2MH
fYev3FXS3on0vfcM1rPlOe+11Gh5RbzgL6VtOyR7160wuoAOHE1tcUEA1lvugibGnf33YjYvQY79
t95raQfP49QJ9X7fDQv034VrDa3ZcMxyzts+7uOCXPRCFHGfPFgT8IRQZLHhaS5DL/4GwfC/h8jr
PVcafbHUluFZ3rf5dTfoVcMNzvTmYrqw/vOBBrt8bXt2IehE8hGLx6staO+LFXEosYKDH3uyBeqO
LpY5Bt4Eg7/OctV1dkHTdgW/exAr54o4X09v1u0x+t2EHIKg238zVvQTkbt5Ni7DcVSU6aF0APN8
tzGKbQTVpmOJeWf99kw4XrvsHDWCKE9XzJ69Wq1QCiFkT7bdOHk2dokxoaLO1AQ53zwjptypP5xQ
9xxMxt09OUTHwGxZe/G6IMdVmnBu1bdr7O30tYICTO/4sPDzH8Q0npE/0ZpHYmVLxw+9HaH//Hf/
MsXizvRqejzh0erEQQ+U/YLtGzdER+CJ+SDuu0+dIkGYIkIufAzvoxeOFczyEtC919V3aPhdOls/
kaDs8c8mReaojVvipLU7j6Rjyp3627JmW2wc0i7cDBLNDiT4AUN878MIsJe+5pB3HgU/VYlmhh90
o72/79QPEdZ7GPFhaUWE6rNaq4cd6FUCEJ6+v8NsLWtdrT4fBAw3OryW3iJLoUVBGQEikoJzz4bD
4mrj5+W5IanoJCwUJMB9ViO8oYQexlp75dBiI067qIe0GVri6I3zAw4xbnT9Qlz1hEAl9wzNoBDM
ovKNtT7Qm2yYL33y4CthSOubgYGCGg+w6pEvb3ZeZ4p7ppHwVO9HZfUe5WekBqda3pVoafdGFDAl
hS5fwCErID+lpBX7wzEd0vy7AVV3fgNmvsmfrnsyBIzBWlQpAeKIYnKhP0iKxfCGW7X1PuHTsdD7
NYqN2OZWO1i20vE72v3My/82YnGLrU54b+N/bK2cC8C33uOph1J2o2tpgM0HlGicS30QhhTnXXoL
fzbqDVOsu0FaAhyypAmXeX2UcWg7dRHKksRR2l8q6w8nB94ZDraOlupIaeBwei9bA43IFI/COe8v
eg0gMzkFgIB0NKPcWZMcSAmkjdtTTMFm3DhlNURbk8uCXtWmtPE8N768FWMRrAzxy+d83qmV/YaP
E8ycBXclMCiJNO9Q1yp5COAVNLml13t5mTwqKYCmUHAW8JCGZ+bwwvc/DdvabZ2vgYtO9b+BxML/
ncsniAr/ometAkQShTAw8YsVSyrTPiuB7GvjLN70jvTGcWMu28H2AigskxS6XlwXUerPy682UqGa
ZZTfc/pJBBFbiXhcqisPbN8P6Qnn3q59Qz1PD7dJLVDRSuAaF24JVxOsBv5/kQbQWcY7KW/NKD6V
/6mTEuTPMQL8q9xDlU3fVjUS4ZIIcoK/PargQcgpP/m4m9wzbjV9/6ks0yeCV9cvcBx6HxKEwrtm
zJGAh6C23crjH1ioFaezYUfoiax2a/d/WEhotQaY1WqsTnV9P2UsWYaTMvT+YIAkekSAuRFy6Dia
9UCTePh62ehmULA0dUG7sHRKmVYsMz31zKCwD9sRaybCUs9+v7i2L80Y9rSMeCVKeDlhpwz2lg06
PWaWQIM0GFLGNYOmlC6R3TRKVjHhvBGsQTlk0HOhevREtgxiL2ZSNq8uhsmMWEyYi2Y50zpXXRqe
3rSdHFcFKXYVLHFgR0FeFFPocD3U3acBX8FjQJHmbt2drXaX9ZefzOBcXDeCMD0MlczZygkl6C+e
KOK2CCDz6dFGUlY0it1O7OiN87fsaZfMjFY8ntlAsvEz43cppMQLCvAu6sfRXbd9hlC9XeBq+uzZ
FIEXi83UXOloP9gnsTx3ftLxzG+y5kFaVzcN4eQRPJaM0NcD9GgFuWVzDQpNnKXboV2nhYufIv2q
mH89biUlYty2XezO6zqArH6oNae1p5f5QbXAsn+fSeLcplt9qy/WvfcY5+YFIn5Ru6H/HuMdieBI
/HarQlNEoS5dKM1fxiCHygvvCKibQlr9wFYaGUxUdPJtLtbG5C68ChbHHw1kAkNhLskhOQU3eqkw
8Syeyt6hbAGhWIrAJsWSxiRuek8/ocVWfxloMmsmttGYwKaHm02mZWJcW99C3tNzpHCZzzKZWWEC
JBHMX0bzQjOuRgniizmIPNu4vawBWZloX7lniaj8ApsqfVkyU/C9MeWAwq62qXe8ntzQfwh+SKkt
l+6WP7NufYw8xFh/oIPWhjbo27FYSxSkxeIyIEo5l0IJgTPi1CQbiToqR728rf9Y2EeMH4LRHyHv
uXoQmr1qWOfaNljRhzrVVGd5aUBR+Ytg/JAfyInMFvpw1SXB/benUZoETFtQXiCmbq88qKptDb+g
9QR8U+r3CLQ6E7J59kgPrZ+gFjZ54tAGC/8UJlZrtVpBUKszejLRMqQ/PJPAX5dzzyehpe/gOit5
jiXwP83PzEz++Fi/ra/pC82EkYCI3Go0RWYlbxuDQRclZItgFSuALUwXi1WStdhm1XVyw8GS0WYw
YunSiJONg0vfCYyWAwiDzpWN35+Tp4/7FmziDqM7rDyUd72FDr5q7qo2f0CkCUC+A1ESGKb/SHWL
MLgRZwxrQ6HLT0+3Yd8m4ZeZoCEyzgX7KQWT6vyZJ3dnp+xOvQUBdLfJW6duVzzO9Y1Q4q9Vn88h
wgSKijN0Llz5MZv8AdoGdJ6zgYp0sn/Tj1am/HfekAt7BKCtrYYXaC1ii12U/X+r86m0t4shPPAe
ck6OpFz+0MMdcf9WKwvkhujkCQD44E9BUBd1wdyF9J6C8xuVeVyWnVlvmCYTYjgID2U0OdthL5b6
AjL1MPr2ixm7tcsBfT/mwZP/0Ki1c4N5lk1W96RnLubE+llP4ekQF19UJcdw3SBxMPJctR/pu1YR
NZwDBA1M61VZwcTuVZbjXxvQjG9+m1BpvKVpxtSwEeGkqXy2k/MmBGvGTu3GJDvBaPcHRbF+8Sn3
+DY4WGNpYqU/WWbkcSk4LB8/GVgiC5pfCWSKeFFy2KYr5W5dMS6ccPxD4HFuyOTvfHNn5G9W2xaK
s3LB7A74r9YS56CofgicMNbufRn9GDhYU0u2xi+bzFEBqT8TuZWSICCqukThbtZmYoav0tcL2p8E
XneWvgwiHOSVePmlBJpXI2KXwj/P0cFCJp5H6aTNB/8ysqPNEdkmYP5+qpPaXc4d+ZOW3kwuhpdK
aTZs1SIdfLo+GGOAIciqEXIiUGvPVyF8XfN9fEr/pL1xvZDQRX6W32W5Pb13UEPXSZHLXSdAImkh
LizKdU4CDRYkc9DD1wV+8uRztFjx84PY7yo3ojHVolyBbdEqtH+IRsvk1PEVaZnuxAxD2cYCES5k
6FJUu0fh8RGckda0AT2JReGmBkMZHYFeH7ZjiiZ/cW8eKGZWVFG3IKu3RUYgrUZ3Hg0u1xrNS6B9
MvooQ+Vlw5hd+w494SQ5Nzwo+f/hf5OsfFmbbWBpyBKkc+z1o70B8jifp9zawp2Bt6uRoCLKLkiA
nwpehS9MzYTJ7Yc/PWCmq5Y4OuffT/UtWxVc0QYhcF7guV8a2w76wOThOH77u78RK0Xtn7o7cUZz
+OssIi0RXBxYiWv3QQT60UqyXGrYcmTRU+5tKH2Ze3arFZWx6PlwKdO+8/1JhpuhddTM3FFjQq9g
k0oWI1nlBypgirdfWDTY0bfi7dAh04YjrUKUcJMmMsNnr98gxcikO/ezhUS43IUqnRJ4ebv3w25Y
d3lBg8X9aMZc0DeQjdt/6CWOPVY8Wza/4/x+/VaagfqLwoWoVS7Uak4gO2ZStWCRFN12uQ1wTXbH
/LqDC3I7ozqYipuJZTd5VlPb7c1Ottm288nqDZWtopvZ99FEdoCfmxZEmYDDkjPwjM2i5Pz6GbWE
7gLelIYWG4Wk0n7tPAmOY66oVwTxJ51/POdIPM8zE4KZoBje56Ki9aMXZBk67m8A1j9u8CVjMY9W
9h5O0cGsPi0fayv948bb7Uy+pcSRTB/fEvKAw9epK2tgz5NA3bcShqcqwG9ZMtjDZ1HRQHJib43K
RD7VzV20R30kAZZx/f47QAyOBRdRKWfQJsGnTYgIm9tVaEMbbhAFWchHNRAjh3Ie/73vJo+ZukZW
Rm44vjHnTgFwztHdq2DFS0VSMYRDvbXdOTX26j6QPYYV51s8emaxkMlWi6jTe1mc5fmVXMCyQMtN
YyCuW0sG4HDk/wxECXXiuG14qhij3SYKUOKqOnFn8duMDN7FzUc2KsBdkRI7XIkzpzm0Ci5eTIOx
Fj8B6OLONxlzh/8S4K0cR+mYm93wLe2s5tSeOQvrmpE0t/B5frFDIrZ92wiYlyL4PzXEZvPMqv/B
WXHJJtHrUgwGEUKDDDem1D2y9rArPQZ963JcPr8s/YENuZ1Jlitv0iSibcDXJn+X1t1q/lz4/z5i
aMtvgdkIPZhX5rnm2O7Z1Jzk0tqYD0EAr78FAQEHNkb2MEMbIBn7+qfubwO3/+1IrnWiRrXBt6vO
4jRH0Zih98pI4eVEKJfXhMXNkPt/r3/V65O2H0jmbHK7zbFdV/y/VYuvGn4kVsTxhT+clQ1kCUNf
cAmE9Cgd7iEpSkYwU18tcvkRwpeBcWGjIYiiXLLRk3rRwPTY8OKEo7Uy6JBJT8QtfOI13g6DVNI9
nTFunyyGimWQNAtF/WQ5J96JX4vO6gjJcDqkyWIbj1D8aiyjPOjYT2J+T0zLIRSX2Cj2VO/QCzz5
U5jQ25tWpeG/kDYH1ESdlRmB2Rb8Z9u/LqgSXJnkLPgZPX66OEiD5/ZFruO5xZdLm/3YcJzgJSDg
kR+0WN3QKwsqTcPtcTpM/4NmFRDLX4sqM87LxTozXGOepPY4kYnVXBE0ehwTyh0GgFX1PkTv8dm0
EkAst0YmhgD1qE/RwLxqZ6oUuM1kFkq6ryaZThyN+IY4fDjTlKRxw03vbsdZqAxmZJu/nDW0d3Re
wzKhBAKnDOFUWf1przRWMijaJ3XadObkcP1qoMruvu7L1x34sVEP4nNTgkcBkj2WHXWS3emjveSn
fkAKEoYlG/79U5UEkIkisBzuPy6gH9u0V8lVQ9QUNRqVYDjux1zP69ldEJf7AZcKyoHWU5Ca8T6J
wGPjTyhEljtapQR/2q2+mDc3XutjaV1Si6euivK78+jsz/amiReL4K8r067R+dsqaMIRa+vsnaI6
Xl6t1U5SGevNS4QXAW0LUucQ69Q4rCSAPr473zWSQt0g161PfWSr7bHjUS4uSklfsBODXt2DvUPV
QW11X/n0bYXGsYEJCSon1HrndG2mW9h6PaZR1kKE2nk461kxte3vFZhOJjlDGa4luIOyAwLyvRG9
KhYLtvk8c7IpeHjvoPH/W7ILrlSVgvxlTIz+Y9ZsU8XmcfZlLU17iKH7QrmERUYICM4BBn+DaHwz
IDKgUwNjJkIoNF+ca8dD0V9n1N2s5Vi79/rEkpKYOTJFgrWgZZa7ull22duV6xZplj+fXd6mlql2
u6/41/1mEf3AWhBNGEkjOxHB8mjeoHf51i9mrqDcTRvOVoYUBoQrrzufODGY1j6VTxidbvNZieH2
SsW+V2Nv4z1kYy+XX9Wvc0/5cdiBj5uOiiFtu4OcLl+gYVEIKgJ7OrDVa/u10wUGsIJQZhJwAN6U
p9PPOIYd2eaOMXC0sEXeBPSQkS+8WaQW2aP7K49QsUDZ10Nc4TjY8TYEnGMgZelFZXJMrFPnGpDY
onWmA9sKTXPrkkhvPO5KyNcMLskAwjKWCE0aFdEJAv7dM028RImr9bBMWqSqDl7u4d79s1QZrYo/
uvmivcAomk7ddTL9KicFjxzEDQKZq0pI+sbuWOlavHN7HUpAoTiKRR/n8mkYMg6Xk54kBn3EsYR8
gEWnTlKJKNtM5e0gpzxNH2kdM8ExikjMYOC5AzFgWuZgK2KqvP9nRRYEn9DnvLwApHbFxqaVNZkz
3NreUoxKRHBMAunRt76MpItVy+P9eJSALUK9sBJo0OpKzDdk/2lm3Aim4WD/wEsKBe6U7PQYL5aG
98Gyd/Y7taojW6VmUSg6MIF1Q78M3e9QfMZOfZDOrtZPDGl963wFhxJ7wCAPyAhOmpwTo2hXfOgt
gMfwWHU7RxFf/tSyeN9MkdgsElcuIcnOWte1UecHmd6U3GrlL16ceRXgWU+73rFx4PZxw1vtHA21
woOmvZlaO5Sg8uxLVmjjZXPPimxXIgSPuSh+13CGoW/mw7v1ineK4f0CGJvG48dyLp9r8IeVC98c
TFG4O3g6NHj2Z8n/hNWi3TTkIzVPq1RqHc7/fWKPqaSHclya+M9evPB2TuXDrWIvNUQQIIHhWnDz
TMn5vBt5rOAKUpNQjbCL+ocwQHpLCdmuQPC3qsADx4qF3RYZ7sBpRrifgGCyQmwpHOcs1bpDo1yE
tSip8QBMWbnAyDPZ1UWqMWP+YEdWFt650tKRoiY75bGK8bMCdoDDr+CSGyeHZbAB/UROXQUBVZ/q
qDccXpekWEqVHjUEvcVfDYbdt0P9TaBLdEpFa+Td7ruHtPTXaVyw/zkCbR7IvkqJla9wVhd57Vja
ShDPqua0M1ZmPzigzFzlu7a8p40tUPGCTavdb+pRXDwU4vsQOmpMId5Muk4DESeJq+iURrfxR4Nd
0XgTGtxCZwWuMYXs+/khA8a+q5QO9sjqORaCa2iuCA9dEZ8jni+6VTFIwRBpQaTVD/uTgByfD7Qg
YVXcUU2NiBbGCqPKHBafSqnrUJHr0TR/sFO3uyhWDhYvymtj5WuxrRDSt8kzgGf7Jpd0eteMJDRE
dB8WJGMC1tsBY0zUPlqGuEzWbHstMxF+KOKIje3hc3RhJrUSbp5dwQc/4qWHoyFIh8uCDSzgIbmR
NFDw0T9AMqOrwWuXJ0jGgxu6WexPGZ7zdC39JbdciFH1AmQAQG88kI6MokLYElT9umS1lp7QGWU8
IS7RW91qx1pg6DgxxxPuWwOsX6W+pFCQ5YfGishxgbocnsbjuf0yDeQEhpoB1vHEyrWzk5x7PEsX
CDnFpY6YY+Fq3tfELnQu8J0eDNj1OMwNYnKcJNzIIeozRrRON/t5JAsyFQxWfIDaWC9NSaagMF41
yFU58+UFl0cV5BwYSLWNoj2Ijg0rbtQfDabhXnk7IsmtevWZUJkrXwF2CbhFcxkyhcaXyDnK0zrq
yon3RRC0sGLUOZYXTtjKadSYkpJS+YcC+SeGyWHoGu5eFN8gPphv1tLwG9YFFeGuZvU7Cbnk4K52
StE1I9XhfgYRo7v/qd/aD9wX3PU5RSdY7cHpWHnm2xNzJP/j1V1OK7jfw2jokl7nn0oSWgQz4qV8
ggVjt78tX8KNFUZjbivs/8SdJsO8tQgcFmBeRGf9gerVmqSS9hTUuMTVviUcmkXxl8VwNaEZnXBY
6RM7sDBUHsGJ3ga0/xKuPFs89FVySi83n2/wZCh+30CbbL0BxtaHjG1TlsinEU0YNz6PovhoiGYv
IzTIwYhBLfXcWqO6gaDsY4XKxx2qYc3hHAkgQNbuPwAv0M2u5E9e4/Aali/m188V5xjTatrfNpoA
lFFT0AeL5lNInkegeWUqeumLn5nSv7LVbT+0f0lZCb5xu+MDD23MdWbNRiJZoVmApij+OPvcL+pS
EYySyRw+5qfsia1Qtt+sGFJ8fPrjFGfV9yFhgihIcktqKlCqUQHQPdnskujncUKHAYAPO5JMmT88
GwulQpNoMhYO/lQOizw0W7FZHAUG1Pydscmo0l3P4BYYcIhaNxN9T5M0k7odSm3YsF8PAK6PO2sn
uqOofLXl6Dl8B8+EY5dLRg37AXVd8b32zc8+kb7Ed8f9xnCpm3GZZXu44UMm5EmehfVEj8lKEAA/
0j6WWtVBTuCpCwfP69hMyFuU58v/eWz2Gau7QdWOQ9Lf/Uix+GGSrUwsSHXlCcGei52fpajLQEUA
laVfIjLvE24d6hO9lCSbfxZIJpu2H+y6r5AW1jUfwEBuHQEYF508YRLaWqHJzyr6MtZJxyMhv3Kk
iZBX2SjXuUP9KwGGlzualrs64I8B6FLMWliBaCGbDzsxQ5eBmUWgMOL9J58Jk5DAXGKogGe18QhA
96LgGFZQjXX5aHGU2daCwrHIzj8lyvKE7s/pLPb5T7IVSU2iwI2IXzul3NiAextCy6L5iu0uuRgf
hwU4stQtjsLG+ZJm7Mt6SvlyqpEpKsXGdNT9H7fYOBvCuas6UQLK1yNxfkWqpT/ELRekOYvQF/UH
W+1+a59n621p0VBDnSqArTkzb+NJK15UFPhuOpoKgANgjAn0uSiirGoLi0AbECM/bWKdfEJps/8s
GFSbFjQZ3zs0gff4GlUF0dyklIzSPvJJlxjRFa+joxPllEcxj0LdPSXfxBbRkLqVfilgcirsBBjr
ubdwIDDqNiS5kJxmtYDBSJ2MZesbL0U6eMgYXLQFS+fiSrpt/W3Ecbt1uFk66aEI6Pd6UKlqETub
vDRKfoFw1j/lKxSqhVTcKUA1iZyKgil45Kc3wte4lpFldkcW/9/rC/iSylI5sSRT/J8eiM0N4ta1
8JjJoIiqZ3ZLUenIlaE4eUdtimfR/ML64PJFOQ6ocO+FZLWmtjQV3fQmcMhW9wdPjidQ+MoRYl37
a+B7iFwi+1lUfB2HkY2L9z1G/gHCuJ/TPVIWKwJ4eC7s/3s9wV7DReqNKaPoGmGXOYfFjDm0tkwB
+fO5t/L5kLx6M85MGuej/G3SuChEMNNixIp+XwTB0JSuqGOMPAJB8IILCKYDraqC7Svx03e+vb0X
zIUbtTAxm65UDVcCuETIHESVbDswKj38UZ5IlGGh1jAdbYu0mkVtMS10fDoepp74wRRUI+AsdKRx
otnbZKae/fhBk+imzBxziFypwzehr44lnfXpjV1IfpbS67woaTeutA2EgoH3tv1Doz9YV+ZuPpb8
QXHOHuwjf+B2dUcdIR6lcbz0rJU+0lWyKkfWN+5ObEX+kVjfO/abh/q1TH8FxOCBuYecyJ/CnLut
vGrnX40fU15WhtdSzEUVWClSJuoeeXQFKtFCtCvp4skyQgOtjMXgLteeh/wt+vw1WaKLV0F4E15h
FBK1k5xQ4/P1SSnBkrbQkyATSkZT5DJSv4zqnHQTvI6wC6qYbeE7qpBN1f0vXLIB91pZfuknmMJO
E164Zu66+/HWbnGVX522/NQ0l3JzAO2XN4Ytl0LIYHEhRnJMBG4CWPqZNm2qgARrbaSr+W5p5mI9
Guq3coBViFeWZHjQxqLL9cvzzI1TlE+bQqTQMO6W6cL/++uF23bWJKewzKMCHHbLqYWmhc58kuM0
HJ0xfESBzzQiynhcb44l/qa9Y1sWh7y7lsDoKUUK9axYIx6A3YK8sH65Jhpvh3ujv7A+13rAoaf8
4yCr133uAtHq+eyoc+6CXzDmyQPu1wDtIJ/RFLMh29hCR+PcBalsmuq7VAh7DDb3Z7MHlKV0v6j6
JJIsB9cZlVmdHwhC/LWBLEV4RXc2BU9ufgSBdtfOsNzYVlcg8GLYaYeIGt1R+jcfa5mb64U//A8m
syf7foljN2FjIaOWnXrEoWNyFFCVgM7tj4MM1uAXXTicJh0Q4f01D+JZlXd1y0HbGWbcBOsn+vi+
hY8X1DnUF+Ou8v9Qfpy8h/wfeIO885HgPRVQR/q0QglCmE2gSb40RB9YialHGg2qG8iGsX2Thk1A
fUWjZux1Rml0OHjdV4oopaNmghcTh9RdnO423II+Fu0iab7O3/1vl6wEbWmXKrAAT3raHk65cNi8
teRC8qu7hGglT7+IlYdpgcjZbOaMA/rl4eaxnXo7ErGvu/ly1fvgSW30x8PlKDsmV8Bu3q+48PpU
VaFAKw8T3SgtAZR/mIABl46TEng6d4xvg8CG8V+WgHiGRHo8Tv3WKdEv3y5E7cxQhNHu5TIm+C4f
VIWB0AjcE2IuZCsqVdidlbzmvbkifj/nviEkEG2k/qU0zh/cO6g1mDNJ0s7bO5X/rTXerr3HHlF+
ZVrQWSgzScCYY30I5qj7OUUtRnMUATiZJXXgew2Utch/wIDQjiM41Q3l+hquybhGnrk5DZXPxral
120tCwN/8P0d/ZpOKFqbQ2EKyF/hCe5+3TuNufYMup1xMiPJsbJr5R2nflGFDyaHIqNiEAZwtuHz
xyaT0F4EpvZaaB/uHV1xJKa5zeA1TlT4SJMapbVdNavngjLwiAPnAO9y21MDeMFxX2YMVvRlbjIC
DY++uYgolYlwVcXku/0G7H//XjOLY7Va9uQntIQi39GToYQLKdJvzpboZG2r0cQxN0lIshYym477
rnW6ogNK0bb797sWIo9i8hI+i0BX5/qfmPXhFxVu8jiOJu6v0XjRzMdFnQNdHGPND0FbSx763Ev6
ERqooJuAkTVDg+25E3O1w4VefBQiUHK4JefJ0HlQtebw/QgHGdHoCx5qP3eCt9aQWAjL45cTRmfi
nscYRZ1ZDzoWqYUQzcGEOxr9C/dTCEYDLIWfTBPcvlv5TE7n6ukroi3ecC9cFiO5loudLbZQ938x
bucx0iWak8YTi35WJQpJAdOpKhKjdj/0spJOSoXAHg2g9ddS5EybpJfvDEAhmZL+S8miXeIBdOeY
zFP12BaTBGI7KvMhQbuFG9NSTE5YyDe8PDbfmzeXx1Fho9FCkJ4Iu6WS1rsaalv/JKAjUh3CZx/C
Ywl1JKq15SZ1VNfQB9oh49Uto/0mt1laPplBtgqe8CGUCm/+aupws9lbmTN9UauYb/CjdR4d3HHP
G6OPXIl1pZ0nhEoSYAVf99gHglZ7hb6K5gTDxHDKiHUjukonjNg8BQa/bBsrdB7h1ABa2VWqu9nX
LRgCE80XzuUnG+0h4fityf/D8NqJNuAUR+aEmkmrCYEWy+kCk4H1+KkWXNW36o8Zrfu2Pcg7F77k
LyZC8Zjr3IQGwRF6G8OXP/LHeLzPaolA/Asg0tJleqRu7dQXYdmbTgPLvjlLBAHTUiBd9qC69Kpc
3MbGczF7cwjbJLsgW5q9KDOxAGqp9cfXx0xTptj/Uz1qCjF8hFqigwgLM8laYd9K+B8W5DBA26vU
6TNXvOQChFSZNb1wyD43sDDkKysv1aUwQoAk8IVulOl+JiiWyWp0jkUWEjRBOJ87Dz8wt6iqVWwK
fsjACnFP0/cpJGRiZMQdUG2BZFGUdbv0yBVVRYy6ng4Upgclc/DpRFZlfmovoK7/pfdRzEvze8us
8hwAEpFRQxrk9af5keOelc/36cDFrjxOhs+MPpBwP5iPeUjnwsZIAwSq3gHw34UzvGJNcUxAadJC
aUBd/Jn7OSWOpGnb5ElG/3NsUGd+6A5RAQgHLnFS7U0VygvbUVOJs2hALRKkbwj3nMgZa2BZi5Fa
ubA8ShGatNONB1TOROyPDxCcVAQzGUh/LUNloQtVkDM/iOaEixNAWg2q+OqmnTZmwFuMhgysuPnA
/WyCpOGkAoudYQHK6ZJ5/MfSaqJDI83+HM1lyHaAJzLjfaVr4n3soVrvd9MXHH3t1IhuQlxDgMSS
0MBg9a4teVSs42qJaqUFR77nkFcsGS7tP2jR8rvxtkLX6TQKbJrnaaRlP3ZKcbFWYFfXCONxyEOy
ipiYkEZ+YzY5wkAhM/89HCJSBBq45C3CowzxkKvVuRxAKmAUoDScw+Oyjmzdoa/SW2fb5KQOa+Wr
RAt7j93bA/EmWwfMcr/FKlNNVVfn/JupRw545NEICwu1G6G/7t5+LtOaAYwXcgOAoQ7NPp4rLQxX
HPZkCdXM1t5Cvfg8XYmo24PHpuQkd+XQRjFJ2wcsMA02mtbjqmpASZsegIZ+yDA15PqItCNXyVI2
f4EsRyCqkJd8H9WHSFKlgWFx874iFgivWaCuWr5CTt/n6Dm9XRkp2as8kA07NaocGrk6x24liJdV
3Ley2y3wmme9xhKXE64EOh/5+Xs7UfOvQmxgkugwt2SfRbaYJgVtscnuCarUI3JsOY2LNSynLezE
ncUomtGb/WJWeyHF2zT/3JQ4HTd7B5faz9+ZOzmWrGvasYHQZpMpJjBcYxm2Zq36DtFJw5DLe4xv
GVyi7xavHMWJRS7hdfC+q3Qhd2LAq4U0rgjq+WYf82hCNWgvnA9SQexmHpCd13UD6QiAw/u3hyUo
a3wiaxXwWidEq1hyF0mRjnqKo2Hb/0l7o9FR1/pR3eUnz45YJZ+ZdCovV3ZVDFNYURYICloj7JUm
vMFznI1QZ0A1iznu5o6FqZfaa9sy3GXNneWNiiXznHSE6oboUgHLuBWP8CJWhZAVVDl8VFiBNwqi
I2P+BiEVjXfVUclbivqDSl+Vo2CvOyDuSIzLLxw+k4qoggN+miGeCe26F7NiJ6fTRuygK1a2vitH
IT2OKu7InWqq14Hpdp/KG+H7be11Qc2bP2BSYMnWPZRzXtm68f5gyoSJJOvEf3cEzYafw9ejLllz
j/+MFtmyBbWlxZAbzjlothSmZLalY7PedZj4AmPiSe/ktjOFRsdzbKfhYUkjnYX7n8XB8LPRUn2q
dFHk1SNxHJTakEX6RL5KdwtVu21jsocXi2fNH7zgxja/acycl8CDGksVmXXablXYBRGTUMj/AWIf
nRlokDXLKaX+NVLVe7QX9FgLD15JGJsqsmjVw67xXYJwOPGKtK2J6NLmSUTUBHIC0pNVivrfxyBY
tDGh7D7DcYKSF+3xw/L1mZOD5IeTfehPqg0cSu6u1zFNKniD8VDu3lRgIpZpgTfbvio2wtOfE38P
Dhtj+72A0D9DOVlQOaw9qbftOKNMxqz/qiVyyCdhByBlFS0xNHBBjUyYktjU2w8pt3rKWgesQ8dB
qbvkk+SOfw2TeHCkUABnqiNtTvkNbhYn8fTm7s2J6bnBWMkdZEY2Y6vuY/ml3XzRNjjVQIxO3KZ8
IA+lF5dkctA6mkdALl7cwmivnRcY70CEtdDJq0oUSSldcWtLfDYkBGj71xRbD0d4T4L0NkMKgUlY
FRJ7h8Nwa8pBX0UaHRuVzB4YNtHNsh8IamTIPtTuKlW/h1I+sOQb4Nt21/1J1fPegBnw36qeMG6Z
zm9Gn3xTg6cy9LTnFC5/drvvSH+QWiEBtDx0WcPQ00c9t8R9t9X0FFIGdKwuDqODme95Xbm9BIbD
RWpUgqAV47LWe84aBHXmHEhyBURfXsHEtVQZo06BVVNxvn0GswP+LNVLaLhVk71ep+NXOjbRCcSP
kYP6hYtv3/z0+ao+G0STuyRmIDG81a04hlsPxAyUlej/IIkMTpypNa0ESVkAQ3tZhIgv9XMUJ5FJ
ZXkPfbNNBSwOJRtN0lm9hcOSQdSsne3WMhhSCn4w3WN5j2nWP7BbcBK4uYHHVtbQt9qsG0hAmKar
jbgef+lcxkeyHeZCCyjK74A3iABLw51iISKg4uKoLSw2AD3gxOUd9/QU0PASnbVNc8WCBU4Zg8FH
oz0uN/3OjUqeH/GUJfK/NlvGUIlSpv8It+83FyZoF6rmui0vUy+sF+oQgRpgGJ1ss7D6FtaunIV/
MD4knIj0ylxfLpkrJ7vEWPefYVm7TbtKA7x77SFyWcHvH70ehBd6f4MDBtrHps/lluwQUbrGUo7j
nwpLUpCTTr6FmE7w507ewZiptMz1LE090+L7G0IbwVTQubuJ4NgAZ0ndE0qlbgGoghxOjnX4+fVv
Klfh0hHoJnfNXnvDlhnUmqQMczA3ytX0Xgf3Cm2GDq01Ri+02/FzvyhDpnKGc1Q1UsFv0eH3n8Pp
15hnyLgRkMAbUAdfNBF+QT7xRAlAJ3ZvTEAhd87aQ0Odo5xZE5ar1ysreavoi+EvYJDsX4luefqe
17hH/1+AfavMwRsOQbrSiAp03rfP0WU97QQrtyy9bcE8FBVqee+qV18eai6clN/QPSV58xBeQ1Ep
/lRyT438j5iQDZLZKJOtT6WMAhAOf7x59A0IZsiYLjZpcOS0jWHZ3o5puSa5J49abH7LDKXJsr0I
IFLFMybLKdtUzWTPZvj4A4NeKewTJPnLv40sOTiyE6ypnib0M+KC4T6zD0aCVXFhALzP0ukmWoLl
SrwCv7+NcC0i4qDQRtpFo+uYKc4cmSoSkxvvY3pL/Q+tSbrexJyQ/qpb03rqHXGVVZo5VXrH6o6v
jglIbpPfGL32XfC9K2xCLNW0XOQAR0nL+V5epcQjnHdRmEd+rhWt6AbenIPcLMbQgNTQTTYqQzsW
j7PC3h1dA5OJU/2vahYjJxOhvNJKATW/sD5PYjH+Au9kEI/ccL+TPXCmK9Xz3J6dJsFwdOf2QnzT
yiKqWO5ev2ULNA5MaKc5QibA3OVVSNcVx/PwcFgno6WSunKowMA+iMgk2vkxQjQ4JlAmxtrNdZgv
7P252mCUwkIUND9WuoMi41oGMzY5yKZ+yocXrQXt2rz2ok3jbnV7lsGvJSZsOZ9PwV/3VJx18PJy
VwiQb6rjcx2cfXYFWO2gJgMpQ3lCLkWP0QFUUZSQCKCLRljKB8FOhIE7lVcz1tB9FzmcRiYycTEK
J/oacL8mMWI+1aNlATLXV4pU4xIKLY/VUqkz6t95NsOSM21uGN0OKo31T2Trv+ONFpKMnuRobRYx
2NaBklyIm1rLcinF+FLLm8bbetDN1kd2XwBfp7B51FcYSBY1SR7JCD97tuOaUZZYgQpxnlWSHXAT
ZPWmFYsQf2eBzeHNM6CSyYrVLmUn9DeYVVi0spINhOJofnhUTG1iw7tkTvuPJMsKnC4pNP4N05Id
U/KujGkj7AUZjMwKajKGO9xTnDABVNmDAOi1LaCuIEcgwE0e/SaPuhUAfRtu77rS/wgoz3p/xj1m
11QxarvfExJRHDWediF1aJBk8UXtYHCxVfh0HJ1egy4H2D5QTx4ulFNov5RX+hTQFfU1/AmJLpNR
Opk1fvMc4eCsMiJNQxD9h5rVqD1Wltsm3e4r1XUFd8WhuCWkgZKwhmj+lCj9GjZhE60Gd7PZAoy1
16bZeyMrbBGpJ6O/J6flGgIi/rUDWN3waPqInWGDIUhFIm0SllIPEwmatqUhjVq35JVl4031YYkL
Ga3nj+BVQMhDYy7n1XtWvNL8p4Gh7yQcJ+wug1dP53vJyklOq9sHQZhB6Eqz4zHhyM8PS+j9488R
ZUtQGEl5W7+yFpVPf875KQSZa201c8yLOkAoKaXmQ322fJyHx3qX2C/WS1VuW9m4SJkh+siKFrG7
q5byYSLwdoClw5zkWHON0K57DoX1+67OolVipCbFXuYIafp1V1/IkvU5Shojf7fVjYU5DhN9VRR3
Ux+Dz84AVbHiShJesuNrFdzhJN1uP6y11n5K0o6M4T6zvAYsQH84ArFoa9dLUrH2ONSYdOgoKf0b
vFmtJ+XS50q/zdr3Nbrx6+FDiKKS0/lbgX0meh84HoUo03EhzjbihpCCzO4GGEcG8alyDwvTps82
zoWUhNLC3Y8Q0JkfEY7QltWSmSGEUgy76HylMzEvCyIcxtMeqYJ2SZj1E9AenLkROFnki+olkWW2
kZPAkwoR1UN6m4jyYK+aXBFIs04ClNibbIdSjDayEhL4QjnvY5y4VE95silIWHqg31us4M9QQaYZ
gwWNwHwR2M49HyUT8OrDqL03nbPm/KcMCfeBUA3mjJJNl7mbdh684B5z0PEms5+z0r4t7hktSmfc
H53VorzqjWQ5NeoLkPAfz1JmiCVOt2b8eQg2RzWMlUhKnylyN0G1NOYWfgilX9US6s75V4/W2kEI
ma4Q42dgWq64LqB36SPGxtQJIMlzrBO2KXc4CUhBMrkhW9/Y5Iz1fDCIQI/IqCC8sq4Tp00CE9n2
b8HWZgLz67zzpawhLD5PzGR8I+Q+/O1u/wAy5uwEEcZTVnWtuJjlx/0ZINi0K3C9tWz5TvtUV7cJ
iZZgQxQVHvkbp9Z3SH4mAid0GOigic8NWf4LVww2vuV/XbyUby6d6AUJYclSCbd20Xe9k+xCvljo
XOE9SkikgYe9+zJDBdBx05fQF7aEKu4gwEQ34pU8BkDh0u5uWpoUVLm86/GdQD5wAMOrrzbIzkwh
XAfE5/R1PNelv6DrAh6sI/s0cDGqTOAAqkMC4vaDryOkw0nhk0/zh7OK25GaOEaLxJa1AKcGZRLg
R36KdKIzgLOxg4DjdgYatLHi4IbPOBTj9f2vO+RcymZPxdXvl1+XcpilZygG27DbN3nZk7+kH3B2
fMfxNLDZY/xJ+iR3AfuoyWFNVxrGf81qwvv922FNU/+b6ZLGcyf0RMQDSqaqryrVd6918o7BpumX
51donZoHCGiMpvMjNRD3+Q79MbjjAb6sRhGp8KC4fGzNH7wAJB9LZsQI5lIr8xkNTrKnFv2OQMfJ
E7kvDfXP0toBj13DPp+zmp8Qy6isyOrv5oHxWc9eDKEPfcz2NGJQGJMKMn5HqYSqff9nDrSDGZ+1
sqaNhkg2yDu8odwklrwMKybHGyJsl6fSnjCK8dfsbMHsdORd23WFyU0prz8MusrQLPGmjPS9He8p
AvlOwpvblEelYwYrChqqQXVe/pw7nR8G1wr0/E13fIbg74vKORwhqxyR6Nz/xFOZA25ai5ywmMZF
XbC4ff7/nk6QYqgFYdi4uOJgWRWALjRKO6+hvMEAGol9jZSNcdw+CI98NsSxuwpJEhF99FE8n51q
HLlTSgT430f7pkAZA224MaprGioZOZ4OymPegiJGM/GunKQ44bwx4Vvom24DIKVGKTStZXGU06iV
GsnuDzgTQttpwlX5VjEB+si+81/DzjuXSA4JfcAGkwDUWGwS5RRA6869yjpxCikCopm7g0uFWLMh
bIgL2YKG6JWLnHA7NzzF/nWCev8OfVe6TGwH0J5ALBtcTlRUHieBacPth0PZhdIyzJ5eP4K9O6Cs
1EdZXRIOG9MWuXifyPfsnsyL3tWwFn6BXyOgKTxxcT9Uu+XZHkptZLRfgwZf7lTVclRoh+prRecC
jhoXhUunnxBSVLR2Iqp+eNmGdsOIK0NGUJV0Ul83uD7moQQaHsrDiYpTXq8M140phB1LE6p8us2D
VvvuDu+41m6gAFi30bbhstFFcviQso0+AbkVv0XceNkO/Rwe5OWCj0KG0zH7bmT6t7ei8CrAftDd
VbRMJ3N/d8lns5ob7Rer5O+mBu91Y3Bnux1Y2oDWw2/7492dnfXVXz1YkhHq3jTSLWEpyZKUz8fM
L5ld7MsNN6nIV4fX6OdmMIZ7KuxhHdTsgFRGZLB1gzD4/X8uTY5cGdjRIYGMhgwl1CCHAH6i5see
jiHDKqtagVK5j1LqlSDIASrFa1cqQtHzKqrITkTUNvpTmPWSQy8jSfYdqtc7QBOluAElPgEMXlsY
MkLuIJXxx2Rcr1vT8LThSCqCHBHK5U7N4L9RT2FqFqoYEO5OM6RjKDmvG5ObR5pVfeZlEblL+4aN
MQWP0L6NzMfnjO2CKrpega5ZIxglMkRhFZep++iRWgdoe96Ph/8hSbEz7NVywrq2+VMBHEb6Py3O
e6I6YGiQwV8sL38N7wzUHh58CrEEfZpyWCTNelg0kXT2KXq7z++4HcFx1OO+htjp3TN7AuLm00Vq
Us6HF8c6Wkizg7oMK9pg5hjs6hD9wh5oam55QUeDIsZbjTol2MRcxwgb9ItP0i0hBGCaDfcNszxg
4P+QsPQzJz1CLwASRKnrZZl8hsOV7vOEyqdTXDVFPd8LzY4OBGm+RKunkeZkMVYpTtYJYZcbgK9V
GlYU69QvlvLFAVWVQbsEVa7J9SRdZH+nrD/te3x6Exv2OtysulpJbqsIKhBD2iJGgbcUIUExeGCV
WLz5u/Zjt+HPoteSf5dtvcgNCdnOLD71YFfeKICJkGWxxmYPpne613LWaARan9UGKK3cDNlIg7LS
CwG5O+s0WCi7oPoiOWRuRpPJU2HsKvpPEfngcCAS4sGQKun9yiSTgp7zNW6sSscQPKfZEeH4n4Gh
z+jI3/zEr/eR5u09en3KarRnxXh9rHnPQErLAvPQ/NXkbpb7IHoWRU5sipaCjhbubQU7mq4ZT703
WsIeGZMF/6A4QYSKLviojwTBMxTlRk3cYCYUiYLeGnIprUYiZjDdOPv5IrucIVdKF+5GzbVREIzO
mGFRw8GwUIU/pSvJc3tNyEABCrDp+MhVJOPyvnLjGX/Ianza6CYfi/vE0kXSCwoN/nm1YJNmu7iV
yHQ4tner5q+Io2T6JovIVOMEp1XN7siImtkyH2w5yyl3TQsZwwrps4889OVs6i1QnAuGArlKDMhH
CdbPFXCTzZgf8LfBx+P7er0VyY7rJa3SHt6Sl/IMqF8nxJavB6uvwUA049wAPLd1tbbZHO6n1ouv
VK4R+3Vb90+AguKHTdIjB2+GScT03fYSvoSfLk14A08yQvPAIDiOh4KaNS8ju2clWF93tsEP1k/m
I99hNeh837mtg0QNgP20Yq51LNX4kXu3vzGLxSQxcpDnVk8798HKHJescw59h7eUOO3A6W4+yut7
i2JlL5A4tl/OqdPNP9yRreDysqO1sn1RgorN9CSy7goDB/WP1mKGspTXQZQ7roqhLTEmbOQVZQBW
rIr5YFxoUXvTOEUsH5AYDLCLfGYIPKtgRreLrOZXRN1cDbvC2l+JEInfdiTMosYp+stehtoEZqvZ
x1lLiFQEjWFNPplj5k1UocRqib8PSwlus4ep/E/q8sTye0SA4qSX9+6QejTm4S5xn/M/6CcsvG5Z
rYVqs4MNGOmLzexYWR+fPF1wOwhb/jD2ICJJi2kCHGpfvHbjDAvXhwZhwivaYcwLgVm0rtIupLU0
9ofHKOIEMabJxIh5QPxGcguuOosHzu/1ebrWYFX20xwXh1Qm21GSAihbEac6GklhDJB432tS2a87
VHzVk5I2r4L7MYsQGvqn+Weaxxi9TqJveEvYPNico5C1U93Nb02LS6+Zmdd6h9LQV3xX4VtBzf5J
D4AdHIJdlDiz15UR9pDqHaYxbqzx247srZ7k3DC+4nPAYOC7kE5zc75TDvy0Wpi7eTAL0fnubfif
NWpwL3+xJE+eG8z2MPPtkhJGDhhtN6LWFyDYRNF41TZTYPsxqLV+UTctqFboArsJGvSV6GvjFzFP
/kkEhkcf0eWeOTE9GgjZXTz4Y+1Rddh8s5cvRI/VJkvOrU2VsaB7S/Q+gsZFvrTNTy9XTWUzXwfr
9uBjXjRw4opyp7Le+NU/5PnLQH4Jkgwlq3jvPNdmOPE9k+z5K1hmnX40a4g5syIcZDQBW01m8vI4
Qh9rPQzoOA+uszsvztH1jPF37qQ/ZPkZyjoTes6+WfIWenc0oAQOpGR5lJ6fAGYX15xCBucEkq+C
aL2NYKRw4A1h2+tM+2yXEm1s3EyC+PVCtglt3m46IMrzrw50mTFb1W0lrnxuFGDcEn1CRQhHucI1
L6p2vNIWSgmSEfAZ514df7XTBQKy8f2557zjIsDIYHIc3j+izQI6oYIYLx2/1gNse0YupZ2d8atS
TXoqaUTBHPWx9+w5wQRQP2PMhJVxjc3qCwL2udNs1qfi+NEsh4NdYAGnDf1X91D7cx7PRxYpqhhz
bjQKRj8mxcNSiPuBVbKXbKfwOhZR5g+z5E9oBID1TtDgjVoaiU58e+LmIckBaA1FhORgswU56pD2
4dHMVGoFpOMHWQQ1QydWl2W/P6L6I+MCFRyoHtY+pSiEi016rmkeuoAbU5r6obNtlRiyCGx+s2Js
LkWSW5RsxDRf20GEHU2AhrnNBD4G7zHYNGvBF2EN6J0s1p7cTuFt6aQ44I7iOWwxlKKkbyNoa2yP
4ZVKejrB2VEDKp2HSPGmfFrJxbajVhUPeKxb8oYF5hQiiTprwppXTJtFbimeCqdMxZ3uvFPOMqNb
AJVJOM/MyP88WdHHZJfDHd2Mtm1VK+bTYw63FJsQy7zEoLfxKBA5U5NVXXSgWeE0NcTLHfZ5sygM
MTFxBnKBXVD0coln+MkuveytfKUh9x1UBixvXVcseelPeHxmAQextJS3rf/29kQ9oTkm9n2EbjUF
pb7oAlSMsJoFnuu/pPK3D9SCcKSVETzdU/OD0ED/cuh1T+S0erRd5yISFJgG7APTvlk3HzvWWz6E
ns1wLwVysh+06wK22wiySsUyshpFZD6NRv7oS7yVUrjvRwkmuwY2ovSOWZmuhzdmEusQOEiACZf+
hlxwkHn1gWHewrFAaQXeZ5O+vUcQ9CsuQKeLtqcY9pJePjPriqkUZSmI4S0AgaMoeVPirF/tvv0H
tCHNC6t2dPa3Dto+kKBuZ+Y63Ma0KNbpqjuJipJWdzH88gqqsMEfKvL3vJ1XAlu9SkfyG37yQgTx
+OfQLHX0QvIQGVLq5Me86NkU1FCqICUFE45I6PJJNQlGahmu0ymnMcYDJ3DIPPzPbhuUvnQ3rrb2
xrFSSL8uim5ZvVsJj2Q+aGXVn6e05L1RHTkU81flA+TXhaTF69dJUImcocxmaAZbVs6C/ilQHpFX
YEuvPp2vMWCHt8dzqe8EF3yBPCO762k9YWS3oEjRk3AwzdJbHLQnFvRlgrOv/Z3HcWOHxjk3E6EW
Od5zlVNZFN/MQp4pmRe+sxaUziiMcxpSQf9nNWIw5+DsJ5qq5MAsDVbLphsjboC9U97dl5Ifpn3a
Lebw4gTKekwGM1UY6YuWBGZ2qRD5XwYMHB4oTyKp9ibK/BY9K3qkPSaP5698qffmJOPjqg6cEYFI
8mYt+T7O3Dl5jmHBgobaxXVW4R/ZSe7qQ7geTTY0K6qoNZOibQdmEaabjweUSzOWEfPjtLVprO7T
xsjdYdkTI1bj5MMIVxP7jXurNkBliSTD9X1klYHkomcomHIfQv0S11lJNAJgcRYnjHkj/AtNGaJy
GLo9FQVpTMjtxOENOD14ixqoo3sDIbE5KRqN7HnuzJZdFPACWbIGyUuhFeOECuvwfrp3ieUgUkes
ycoCk2umVodWIQCTCLsGHplt14C1wAwsyz4ZQRSx9g7uPIT6633eHUf57ASVnN2HjHlAMuuinuiV
pHEm+8g7OH77leZbU53NDm62X8VCsmqdkwK0ZPW/8kpcQFNOGJiijxGlom0Y8w6VJ43rD7ED62WV
7JyZFzOA7PO8r6DT8pH77Q9+Hnw04Poefrbd6wpIPUGp45tF+5X5uJWTHSc1iUW5QEBXA9quGv5P
IRiygyuHn7+wIs2F0y+ZV1aWdQsss6ztWpakijuEu+Q6PE6PYSfz8gYOEtDTEoEFOvsnj6HpfMs2
uM5RGyWc/txe1NlBfMRbbwJh6dT/zrwESwCS3hwxt0VfN9VbFG1dEjWnUddGq7S37Z+qfWOd6E2l
ec6tUXeADQDjGrqb98d5BdgNAyN9lMDmCWXGY5b/JDzxTMTCf56yVfOg9FcCz5lpWa5ZkxBsLb/Y
OgUIYi29V0zhADS8vYbcLJ6mt9BYvtqSKwR+urxBFKz+GWY2kY+PRNCwfGtblKt/sxr4WZ3BPQbA
JVFYHqT7EJw2TmOMOjm0X1vQXxdJrP1g13IuTw3FAFoh5lAA72Q74WMi6HrS9GS982dZED+VKmrW
eeAwAQgkFkW7mm15yK9CRD/5lHuF9u1EOY3pFAvQ34H6bPhE0bxs0smMFWUocNY3IdiW20rdrb3+
iBNsVSuu7IHoSf84G43kG2mokwcNg/RoS4KptAgqRT+sVrQ7Y/LGSK0puMRWl1891Iqgh53SxKUN
MJmnZSQANppnYDop+NGbuzWo52zYivORuXH14inwpWnm8lIzT44tHTYkLyNSr721CJNKalFqMgGB
lruH9ikZSyMK6gMYLzjftzpuvaAJScllVCCKFODMr7r7B9eco73m27LiI3S4HMJPTvPdI0rnH+Yn
Ob8Utst08MdKOiI/jeNGCIblg4cbpRnmu0BKWySwCWbY8BABLpGBneQFWxypJsbz737hxMVhPVTh
JBjZNLX0PwL84fsEBE2XiMvNNMuXCk6SBMZiGe/1YJYVjvBWG4mtLHBRWaPzM8qyqCTCuQa0MMf8
2XNXqKAPrxpHUGVBbG/pXx8dM5ezG3XIMBiVXS1+JM/I0CwkOtgNA9otRO7aJps1e4iV/InkXlJa
mjBCyEk/MDzs+rNrrmmBymvNaet25CXg7o3twgoyqv1vnEz8bb0AAuPC9NINuihfugXYExEkN5b4
GMMK7IuMQwCj6EZ4H1K1LpBfIBm+frzXFQi3tAIBdyNNduvzTkl0dA2udmxy2+50K5NWhQdZk/k2
5yxGNpvFqNpHNWdcJxrntL5RZ20eTaC08b1WlAHX6V2CliRnI5IDLnkl7lhiJ4SCgVOPwK/lkt27
ntlg9uAfAO7oGCn2jzrEcCJTxIQpJWsG9B62pv7Pdz0yn51DkDim0ciJvgzuFyVmINjEdyGlpLkF
bVQsdTnoVnEw3tgAvu5m1oUJu+pkTLyChALXaieZEux0h9p06AYIujja0KWyMNTDcxYg+XnUhFYC
TxdVvW24GiMprUwaJvFF8Hcq5ZmAwx0sujyPhzVJmDju4KPty2v9pCNuJbNjXljppEpd+iUYcIww
toA/Vd0m7snL2XbWPOLXC2nSE5WCKGfmzC/GI/D1MRT5OyxqRZFPLLfQuK4csou50KToMtsokWlE
DFT3RHcQprf9eVPglmFq4R5iazuO7ToZTui0Pj4dh7JnjQNC/Tn+BAEA3eisB1RotJ1YlbcVZ1dR
mJHQyru02znxrYy4v31L6GNTgSd0DA6Wk0x1qykgsfvVokpl0FEJ3gx8VP1bDQ3awZqpAE8MaqA+
WMSUCHmOdvwD+K8KlaoVv8nPfATG08dMqP1+vdBXU1s1xIVGcEhb1Tfh0Rriqly1zr1wQUpy8zTT
P8om1sSVrC+WaVNvjFMkmsYQNuBzRo2ybTCLrNkmYv0CHcvAYmrjJain2gJNrDyp2d9Jbvdv3VEU
S8zCS9Eb1PUD3rf01RAdNuQlDmwKsuGzGNTMC2XqUyPxRkQF2p6OR1Chb0zaDGmH6VBt2C4QbqbK
iS2828Y/17uedp5mTA1/+mwrlWzCj3oAgxQwIWEhu6SMP/FywDdEZfTeSQfDfMJrpM4aB/fgSnb5
kdot0ArC/CHhLYsVjuHOfGs74oPok/zFZgrQTjp91Sq32G9dz6W/vlaiojamHVIDdQqrJt9oZhGp
Y78dMm0erBwpjPQl0vsuAfs92FaMNzlzgL8tDnxZAAdnBc0WHc2THWnTuecvcBBDTxls/qehoDVp
q/DuxLWuzn5jKojMFW2AZksZISnih6gtEepl91ZUQwZik/LPcespboclFUoqosCpaH4yhxvCdZub
zpa5jrJDxamIWnTD+q7aSUbmHqOP7QVTcQsq8IJOwgtr6MPd3QnJESWcwz0IUmW/zdCKtYIyL3qI
CJkUhx7iFxlgBBjgQtKcrtgsPDj1IUXYlfmdJorjJ8XwV63KKJ8RaSLpbkXT0m9+pMCZG+xxkkBR
mXQQ3OYJafeRc4WjuEJGsaKqa3+89NQ3HkmpuNoU7HGhIUC2MUvj8Tq5c4xcNYLcN0bCgc+fdMjy
59amdw6r8RtJWJHMC8M0GgEjvuLgvIP/9RKQ2Pr8g0kRT9KYFnzu9SW5esiZn6qfmXUiYP9pvEnL
jS4Em+PdVEJv8QK3LMTzV8NnWs/u9XyLlFoUaQ1w3aajxxZVu5v2pfM5THt2v3IJ9PzRl4YsrAk0
6zA6hFH4L+GZS13fzOmDW6L0Qt0866rCSZ1NRlP1r9ZOAO2LZHSFEdZJ/5wCLcb1jtwp6GDZ4TWr
PsCipC1NTldpdJSVX1lO3kvN9jmnNMoaFK0bl/W2HILByMQ5vOwYqLQDb9vgLxh/2z8AFUfSehqE
yNeKC2DgmLe/y/hYNntTfZzM8e1+FxsvY2LTg+q1Nx2W1cSEUuLuTnxdK++twxdDZEsFtv6ZJ6or
FS4t6rcgHRCNxKrIALmLrJ8q3WeQsNbHU0tBsxFMSv8t/mM3bgK6s7smbYx4e3GXtfhjkQaG9Zbh
EOfQF430qOcWqzH34B6xDfq6VSSgVTVMLV+BB/DPfR/JpIJhHNc+MnZTkTnrnNXY9pGlGmn5Uoi9
urb0wbMe4qCzyKTHVXqaJmlvRjEpVp3AjTXmjcM47JHbSApjKYvSK0+EX6svJxFjuPZLdzO0azl9
agEm9oVUPwyemvHfgDw4AZ79+Gs76BWgeBEj22FmjI2R8OUM4IOrNk+FJg+SxrRfGsHBelUflt3r
OECQoyPSN1C2BXYVt2mHTAV7k/9Pcmm+Cn+k0XTLbNO5X6/GVX9AE9Vxykh50LP+Jq8BAdsY4CJA
0PbYGXcZUY9HhQiH1uNUFoksf42y9We6tVvK9b+isf+vFbDFpp4bNf0rSkCdFTvJoo/a8igxLk0f
dEFGQ+tqibkoraXMWWgKbdobi2g7jFLPZsjjAw+LQ6IrIaZ2VZMoaNDwMdLeNOM+BqLHFVwIJ1Nf
O5F0ORYuNL+tcVq15K1QT75dNN0xbJhmCGFqXW80tKEFeiNFV5F8igJOKxTtnZIXPyU7rfgyuQ/K
Ps5h+ljET6+b3BICbq32PeSUxM1CHYxC5ZgNdFsI9tmsmbGI559P91PMACIjj1p2I+eeSM0UFahU
mW6kaAmkrrdqqJS095YyY6JxtQSqaxRN8XuIMnI8+owBC07CRu2nRMNGy6X/7I5HbRTWG8bsQLr6
8JSyVmS2qNdtdGDJeVYNXzQpH1i6LHqlzsVK+TpvZc6T2V0NpG6gr8HY6GkI+EgJ93HH0Yl1kpKW
m3ZXnVqp9R4sxJoDvikq7kr/kesCFXzf0JAGcc56ARO10hGY10Ss2Olt+yMp6UHqKga1FNS+pB2T
WjCitSOyKT6FYIE7LDaqNsruHjiifEaBuUx6M1G0YX6JVb+gsj055kcX0O4ew7NTWS8GgCdapgDj
PmXni1DzhIyDL4vcoadz0TAokbw3BXS8gVmk7hmnj3jCeS/0gb0/gH6Y6k+8Fl5ySsI/4zb+0Z69
xShSe3EQTupC135aXUL+bcNfPuYhgDlhTWbuZC2crRWTSfD/2aUv/Y5dwJxWGt4SL1uZNGHBgqSZ
UTX1oISGAsoN80YfTsP/n3fr8VNtd0vf9E3BAi2hGAN61kwB9ugb637lBz4Uvhm8nnu9wzmqxpSE
Es6Ya9+O2PJIZvakbxoiFZoYpRspKq4VgT6xqwNTV+TXQ3jsPWrT8F9kFCZ7oNYXyfv57cXuOKSA
m/4yUqNk04QshycjHIePoTp3ls3OAAG3xmH/I9rTbbO7AAFM7ugp6SifkPgF4cqK6Bdy5vkJMtS6
QksJt/iqotZKWBIIwKWy0ofULLiXPLcRU/gV9Q0YaqKl046pk8Xl5jcnLRRQ5tW1W6nTsCGpLaa8
CWigMLwMswBvFvztHKzVaODAFPuT30JKAZHBvE7zSqP0l6ObX7TbzDNUhRvhhzA3VimnKuqZOF95
hjSLXKZEJ4Ldck8D8gjmGfzrBjF9X9SrICrK482Hp6qB4DbtrbVzjUe19Fh8vdGcYu8HdXkQjn/z
LZfBwG5vs792zroe7RH8Ta5kRpOI1miUtEjuBklPZoIi6ph3TfHlNZS4E/U1Wp6weCKIysLkDSSM
JkGRSkO0YfGip45qONtPHrtm+zaulwiibZvaj92PkaNziHcQqarZ4ncmrCCz+cWIOAjURcXNPppr
5aAaBK8yzFonLjaYfbKgXXrrZCjcnzs8nyqpuGLxS1VasM1KpoQh/CWlt4Ucd/gqa6Qa4nGbg95y
EdEcdF8+gcRZ+Tj+7oIXNAGpsIkLQkNWDPpS9fX1MJtGjrrUaAxY9/4OdtzZeGwj8fVY8d4w+rqW
aEEv8/Q4ZmHTQ9qk+mgLGj0AuCW++TkWp13FAsv4erUFAODqZ6s5kv13zSWrZaeBKo1bMCr8u3Pk
gvAiL9nfTW69BXdWhSlulev5Vd9YnH9qhs+kNES5G8T0W4MGzbiABHkIkz8X4TyaIXejAneke2vZ
UtszmFpssNHOV4MbfIz/b6fQ5tVg8lvTl4eUCoc2EhhNF2mVbb3KsQolVunk9agw8c0KnA+fgH3T
xvOkF95us+vwrgibWxAOWU/LX8SPprR5MKc3DxDJIDVumy6XwB7eTctvQuGlgWep7IUwU71ds0cS
UF+ZCfsnEsY+kAxZs+Zr2Wxl1ZIDIp8QFRTKXCwtpqhBvRFN/V1IqnfCOJOjW9IWztE4j/KvPivr
7eDfaHVRG9yoMxlgstnIH6A/jDS4ZOGMpXyPZYrqcgAte7l3FmU8Uj9aRi0sz6Y41mNPiY+/o/b7
yf6BNqyTiY/m9v1Vuo1IjoTmunBXH3W//ZB4+TYxXl2oeGy6h3YmuZgaJoyEWXSw/Ju2iKbh+Y7H
ZoGv94Wfa+OFfLF3mHmg4bRkWixqBpM64F7kE35FMR4BsM4UxcaEWjuIgyyxdprOK3J9QDtzobKE
GNvwglboxvGBib56LhZ3vriE0gCgWXtxN/CnDak9khCevlzoMTL/L3wwRBQLGQYdFhiXq21lwqNB
y2OZtHuPB+KQmfL3oADmdPjMoOTxdOmKanxO6vuXzaH5U80kKafE5KJ+zbXKtiXucYdxNTmnExhB
DV8R4z0hXQYzTg/JUSePM+nZBZ081+/lz1uQsWOC0DkHjIeu7lTyEKDdp54r00YZ7N0ARC47bPY4
R8HXo7i10xQ3ZHcuu/PkWF+ipUvnkpYztu/2lP2XG1C2MhEqPKBTapO1W/8xnEfepcQ3oBGvgFgw
Q0Jc4j7VpjjdpJ509Cb84Uyuj8XNawQuduPGXU+s4NEdqdHqhFwu8lGAWMYjHGLIqZoTTRgglHa4
oxBn1rjl2OP3I+XDZLa3KHdsO/NenL99uxVlmQ3sfhh53qgqRzHsIV8nQGglfDL8Pob0zg8Wgqhr
xO4Le16MZhO0hRFEbCbvewjLLmrHcC+972fH6NEmihql6Ynil7wXadmWtv7SV+WYYd8Mx6xegDjo
VcN9NJ14tDCfSWtNml1B0J75LBk6/TYkUlLy+jtL7MgNPAcSusaVOi9rRDK/CrUEHxmq4eA8HABA
5Kq/r6sQsKlGoJ8IJcLND0GSgb1Cnl7N5Teb2MXte8UtUgj1ewoa5lRtkkyIDaBR8ofWUwobBi3Y
ebWynFxhE/UCjtOwiP8HIQ2e/fhYD5Mm6mgiMwltFUiBOAvki4WA9PjHQh/1pmN0AIDpUH3NKhdy
EeZgCO7ANRrvUzlE4BRGg6dWHjcqQ1bgC9jjYZXntahHk/957Nm6u7rhi70yXlG3T+3SooFkq18b
ynYUg0czt9snXWjGx5QRkyWyYazgVr4FTO4XUABimq27ezdt+vr+6AHYNeg/j5kvkrwFlpOMVSR0
+rz0ONyUZGqkl/CR4HDwpdeqWhQzDDZ3FLpeVoOinJdlZ3i0M9MuRRicOv6lujZGy2kybgMClcTF
+ERl4nMl/w/5qA+iR+MD9qCeuKJanyPZshZPuG7GiwSf8uz9r4H83w8twuWvwZV0es0fL1WYJj1h
qtyJCsaeF/aQDMYqqic4h+b0RF8zx1xW/kuU7IHAJqPyYR9JYCmfb4nYPhtemHXfU60adSrznqhp
Z5scOzohLj2GYPJkeGQnkN57bOGNCkx9/X77pQ/0yEelS75jlI2ywY/FFPuCnIRSvBG3xqRM5KHA
x0siZ5X9F6tMT3g/yZL8+ZOOPqTWxvT+Sli9Ii9uRFxmtAbPfCO4wiwuMBD2JvFIAgDw2ycvWCvJ
uWnde88CE6OrfKn67Jw6pRvv2oqmAInOE38/Qusi/9OKqH7b/KODdFQKFPcgGaIcH+Qu0/y0c4LB
DGt4Vc+SKge7PPI96/TXNAkO7f9QtosCLTbzkuDx2ZjiqVmrYCi37YRqh8LH4tUyDx4bSnKwpbSd
XOL6PXGZPb/Y4pFjuz+DjHEOnxFqF3XjsGrR0PZ+hxaxmN2LEXqMkSiAi0RWGM9D28h4kT/Wn1bM
WCqBhSKRU2IZOlEBLfcWVksfiOGmMnZcKCWgSoQLWD5kgM1ZQv4P5y8TnnKunfx1HvgtE6lCTH/h
HakbpkKh9QEo8peqIzJdHytv1lSDlXZNxL0LMXmSFMTzvWWzsx7LgV6bkp/Xx2DcktI3X/JvcIWo
ZpHtySE9SqN+Wke26AbYCI+7z/AoHgQowXNFvLXDwpMZ60weBihVv6wwcPGacnQj0mJ3W610gwYA
SChwi52ynxqdOaq39yLfdNxV19dNK+XE9VR7UgOlVQ8HTyhjsPDvkN+F18Q7RTwI/nRPJFjkv6rY
zxJk9Yx1qgpRozXgmh79Rm1jc6f+4dNvZDH8nNuJcoBDDDTYybxsIS+nYcK2S2/ykJFzGdjN9rDr
1nAP7a99Q4v5+6Y68oip89y9/JjDaIGKzj/0gYFZv5wbiL0EQXV87JVqhPWFR0HH042EbnRXUih/
ntSUGpJueryKNMJzHg/4a+Io4vFMjA8y5xHOzaOl+4+uAvjBez6MOuQCngxo+cJIoEC+LkwOmKL8
BasPMDNGX1Evdj1jltFR4XfE97cb97QABnsO2EcGKWaKJqoQ6PqpBMC72tLsI3N6wn6Zu/PJKTmB
uj9U/WGH+v6HRfcrED5Ip0E+6yyv9McvSWR31r5s71EOGxlUpuQf0G6cIqV6c4NFKgwoq4coPICu
G7FM1MVggw1TGZgAaL9z6QozSLPOb58KGL03mhQ1QtrfjWmtjhtcs3Im4rPNqwtHyalb30TzQ+rh
9Qh0PXk1Q2Tq3tODy9fgrmoHa+CWXeEKmmoa25IZuvACtc5Q4NahAfJx0VI5PcnbBU9kYLkDovjM
yApMbDFjJH2AfgiEeMfEGPbtihHJ4Ubyp5Ey/ZQZHQEauQODjZtoD8DVFE0B4fCzlBQzaD46p30v
ohypG7N3VvTAAp4cKK7Ujm7AyLuJRwkffDfTxXNP6a+TWONtHr+koZdRZrAr8evEoj2srpHdt90+
60Kbz9QmJxnUY7z6/hvUGrjYR4ZctzC7v8a3LHQgFIpjVkVUKmfYKuQrWUlwmnty3NssNskg9pki
zL+HZz3mE5Q8gaddfYA0JHTgD65bYfoulFddHp1TTIkGpQ3fU1cPyCfwrlAzjqwlo+TAmikRizPp
qlk+0fgyy/klEfIPYt0LmOFZTwdc1hze1xsTX4HjrwXmyRffJSWafO9eI7TT4lVD080fm5tlk/i2
ITzbHlml7IS8DclgTd4X09cBRYwl/kGFvpg+Z/xCcGY12pwazxdBeGDbE7o8HoyS0VQcth+r/11x
TJKxadao2zhVAJRBkPXdcFwzNBvGsPOQJ/+l9b6kdIxjIvSBNGcYB3y6+tDwOiQRNvVOmeMXnMQC
p21qI5/x/zbWlDOnD3SoPPsWnbglKMsKCzdQ2Moj/s3DVAgQLspeK/D3NUjo8tR0KrRNze/fhncF
lfoH2MtVy3OgxAzFlQFF/mzxvqy+ezYxpvcIWmesx5SmTaLvnfWNHcDuyavcEGQciCFz1Do3jfKb
LWb1wf2Nd4aa5uHi03x3/1V8bRuqXpOaF8OsUWPH+xQlySFgqRu7LBccwZER+G4E785IbzMX9XZR
Jhv5unkeTvA8pI9Qq4bUgIXuizM5TRpkMLygNo6d+WFxmIiYdLBxONC/g64kz9Asg5kjbXy4u4IO
yhkpPfbEVEqhJUIY1uuGRC19mGI6kF51NBLxJPt5i9qB69YfpobIbACi2Eyd+EGYm2v5QR+dgCTU
3bJOtQVMTNkINzIfKwY8omrZ+CF1LrUdNHX0wHa5k+EBUmGQbq/sSJC12H9dxydizqSdF6N/aaLP
2B49iOBrXJhzzPGnN/ChVsEVeBQaiKo2CZrYUGhUOjxQsWKwyitzDt4o4zjjHylpFudg/07wbvnv
43k87GhxaneN8tUySwdrm2sHegzfm6PciAKcAMlhAzH+03vv/WG4NoAvoZBpr+u9D1EMHtQV/nME
EJxLmJudOcZ3m6lyh8/4CZA+bj1HxP8eZeIMr6U3lbTsErpb02G/D7r5NF7e/Wlbxqpj67RblgkX
w9fPD+2PEQm5z15/oy3zsVSTvLZFSHgPjlOTIeZ6JkfBZDzlUOTwlElggwWIVCQlftN9KHR0pkSx
6BTIm6oZIiNEOJxZH/wbbhT5SsNX5RnsQk0w3amqsmH9NIUD5rexnUu44ZqD13jkA4YpDHTCxQZS
kiiV22oG+3fYNrzmOBKdx4QcSby2WNGkkiKUqZyMZzdXIjoj3s3jWco4OMeyfwjjarKFM7iicQjY
YyIIfhyreyB4aX2jhHEjHTqTpjk1nRSiIURIDDrzkm064SyfB6AM76NblWRzbACMN1L6xnnC0MmH
O7ow9Dg4pbDh2DiE40wCPKMOiqhZ1NLJzg1bG7T+alToKJ84ASPy2nkc4OQWIwxivNi0pHetYkh/
bkizY1IsVYCQ+uLCvcnMqchy+nbuQ0Ha6+s9lmJwE5TJ+O3IycR0+KfvDTuOBcovI1YiSqXqGMoA
idk1TBRp/dn49x60WiExe2P5BHEe1dLp0f19Ie54rVjbXH0nVfPDIqFTUx5aV5O0bI0MfgDgXcAo
Ov/NVBWQ45ITOObJcAkL3GgF49cM2TcH78jjIupxssCWIEXhRvPND3C9yuAd2lCVWGs3P04py7r/
Rw73mETMXORzx7JolCnR8HMuBRXux5VACId3NKf95PHMVzPSRO5yV7FIaaJ5tvC2BOXeDaL0zzge
flaj1VcruFPJkqDe5lw6S9MnyJjLSr4/ru7rO23tWN8AHJZ6tKuAo1ZkRxcBcql2lNM6EE8AgPeb
ze6RzUZde2O7/CcUihpFXKqHH1rWqZvi465PJsjJvG95pz0YNTOvpXuLJQT7jYCSWflLgQbG3uxc
tA6xlHJToKuMCn4rAHbbHfWbMv3pRvkp5fHJxO9YJ/FWo7XblLFENqNeAlD22iWcli6/d3np1us/
BT1FRFOI0ecWcNoXgoKPVqpWX0Yf++9CuSmSWBwOI0ZIDBn1bZ0Q3aCukT9GAsd1wUp8vwRqOEFm
bT61wLgsiJldGaox5vSnDFh+d/MgHpBLd+JOn686zh5D7tMyrW1xqvim6AN/llkUtykFfXzgCxmf
RJ+g+ax1IW6p/AhPt/gfSeGjE/A10FESfL7T26HfeI4DR51nIjzICrTzprIYgDu4O23020BvAtEp
zsFe+TYREFPTOGrwZRwZDNITayIDnbfk32uTOxnD8H18nuTlC2lyWRLoyYhYyyy23aXyl1gpZa2g
9HhqYpLsz/kiBT39cFFNcxGQUK8HOJTL0hhRSP34YDpDuxIEWeCUKjggfujKgWy8FvlKANH32AKL
Fc3wIFZ0pNIKoj5EkP4F+LE764+8pKDfS8h5rh7t4KY+Vhn5d3dUdzP/VcnUEbCedDfos0IpQibO
8+jKpoltHxOHIdu6uJYsa1s6VU/E11NUZHV5H256YhBo3Jv48JshCiSQg04xTR8otavloRwHt9gY
v7ewzekFnjsMSAGa3RxmCSJhEKrnU4olLbNQxxonbNk92+1Vv3cYq8sc62ydSVAg0Jf6HiFR/ly2
I9vwd1FPMGuJFKaMLjN/dNVKGVRN/J7/Vy0tD7lDe3WppDj219eqccWxRTvQlxjxxCS0I5PqzOwK
KFpd9BVBO9PUxu4+sZMcVpBnG2qXnrZxvG+s7DGlhIt+OiSrDi43n0BMd4padke9rnVX6+BhtXpQ
90quDm6hfi+o7dDLCX4Hu6QUqKcvX7D9cQ+Y9r0sH9gtKOKZwaES2Sd4CusCGqqz9+gYsXlCTBQ6
On8mxFdJxcG95OZ6gnZ9DrItMZFmmdPjc9PT1av+BBo7spIj4WuhZRkg5cLYIPx+kZ8HKPz/mHXF
w/omgOLTTzXLi0pdWjp9JJ6XZH7+TAhWCWCxhiZNiefvoG4lun5L4fmBbeM11Lhb5W2N/Wb84706
gRXHIIxEv2+vcNm7//FXWLs9tBtjXLRipks94OCcTDOJi7X9cS6oRflUlcHKnfj9oVdlpvouLBWs
kJeg9dVXk6r47Ge67yd79K1M3dnM3MyTRyvIJDUJAZj1HaEGBzjaTGHi6WtitYMycddRY9XBVlqn
ANSJf5pcbJgVgiIXMyZ01SaJeQqWvKxkd5hUGJcWYodYjkF+SACTHggRbFkMxw6tczUJZK3KuMPY
mFGQkaoixZrOt2iYe18+fZQ2zV1ycmBC8kiSKJCVPtPnHGt9k05hkSHBzxXjyHVl6oG9fc9ZMR7j
ujoctHlxpXyGat6gQpbdvFpu+WQsHi8sQ+4rWgLB77yaqDipDF7cRFxnd/BDZ4OqMTc23tFCdoMk
tzpKn9DvPBQ9BOhba7CgAvf5JfPJg6qzMaUBdxHzFRXkCke/5y2BTUxnqzZnsHqbOVAtyzayLGAn
aFhhiJDopK8PE4RycW62ND/ut6R6C9J6YevG1W3QxPIUbIok1iiMiQTaPQqFqtAs7l344Cw5wMbL
sHAkDTI2T2E3kxzyA9rWGKfVtQ6LmTpgJpuAPJvkQ0NBSKvFgpyJ/3J0ndAI0J59hzDC+zqtb4xL
XZCXQF8iBzDm82aP3m8LHgxBoyPO/gRAb8QP5bOPLYAzOQ/7Rc2U3Fl4vz79epD85cxjXWJkzQPK
mTKnALlyBXhY1pBqXoEEuSO3+qci4Ygd/8dyb286LXK6kOjvbjISn63OgyKHzAt3HqRqMjSllPeW
+2gd1ewemDmF4x0sXRcWOZGDgiaFhCWMZ/lETeZZr5ZgKRV4FpvGNIyoxcuxXrWJ3Uj6i1Y2XjVE
zG4qlDIMYmdVt68/3+WLkF7OkZZBaqPZZjXhJmEvCjti0EOy4rB9sdAEkFwsXm/szr31F+ihqQmg
KYF016dLuDFccQsreJQ7hL+qHEkdHJZJzgT+sLxZOzAyJToCxC9Yw5DQgcEF1jAEU2hSWfC6ddHK
Lzjwuv5/iFqTujEjSES45Ph4gIFlDixHVfVUqMMDAmSzrBqGIpSUPYuMGyp59d/XfbLkge7/v0wz
v2bJfdMqizSEI3VifFC/8oxFimUG+eb9cTBFlScVqH/v5ugX2H0sYjG7HultWYKkEuzs+sGfnpFL
U3g9J0y0NIjjoqODk7brXbk/BRQNbVSKMVZUr6uoaHxUhghgORGVOgpkFA3ptImgPUJlJL2n1VkD
AIuzyUp8XSJv69a7xEfhaR59+cN6BNkyQaOBhr9za1jmslkEUbd/tT4vgFv4ieFN0fXgO0gonBVR
m5Fe41HFwRO1JUA6VHxLDIN4ghi0BxnraJJtNvIzDGmi6j/f9G2QO+/fQII3f7UoUF76SHm/CMMh
Kf3fEHr82Wmuel9pin1XOy86wYnXO1NSvoZHsz5s1oZhvgATS7YFWihzLu1NDiRMNISqX98arcDa
TxIJ8IbR5s6zY4edc+5z0rbnChJXupgKSh9lYvgVUmFRkxyFl3GnUXCxbBZaMg+Yw5QGSyqZpAql
ZOSoNJ160+Z+75zDZKBW51skJJopVq9PvMenEJSL2ULW5J0UesWIi7PUKUqYMB7JOau+zIEHhre0
JFMAm6yWgGEr6aK/zDsQ0XP+egpQbhugWJ5tFJn5i1d8WJhGjvCp1vnpXeujAf6OK1QiiPl5tc0U
lWsiXRsjrHF7S+cdyxYgL1GZ6erHX5wDAGjc+bj7e5FRAuRfHWMurzHtW93xwSw4t09DzyNdaXHm
1VnOvI1MrDD5L95ZQb/wyoQY5ExmAjvfFQiKzCtawRQKBwSp7u7DCwEcb7hNfiRbWKmwVXoIlQYj
B1FReXDKSCwjWe4bw4N2xJoK2y5FYhZahF6ow6tg54QvLaMdAlOXjCzZOOSu2AycVmMG94a7b/7e
Wd9HIg/ooeXV6M5eANhdao7lY7MguGMhAj41VuCjlkIF3kSVYUrTyr2atq1W88gMw/6fAAsHd7/N
YcTatJ6u4dH/Gu0MrTiYars9gnGLKu0tEd2YlUsxgufIqwccP+QySu8sEiS4brXL4zrSjz9MmnXW
pp5eLbudjFi+K7O4IBtNI9juxm/zQSVi9FnztFwZYxz74tYP0MOPE6SC19+k6CVP3DUlISR/NYHG
uJHYPes2G1gFj4RMNWLQq3t4lariTdM50nQ2LS68vb+TEM8mqqDUQ2DcCe+pHP5WqBWl36VMY+dc
FiliIzZd/9lWpvd1qjmpXSYYcMp1+IwcIZeXPIxGjIJfmjIekDO+6IpxqON1wGV7cuMw9rVEK8Eh
aliu+PWUqyzOGvM/c7O0K6d0ACVC//Qw4GTjdneBqOHbEYs5GakYIR0VNlu9ZuSum5hSOrzqNMjj
0md9ZlJqzgaXWIggywbmnU4NVLkmqjvuflYY+OOAgLIrCZBP4+YUNluu61GXbnZEmsklzKUcPgZ+
EowhFYCw4J3xGXhw0MdStFxcA02B2WgVnp34zRJgQOKNN6LqeWu30opbmShT2Xw6QWV/n3t8HYoU
jLSNBa7vb2X0NB0cenWgkeRUFQqbFhTMyJa3dm0WBbW4ejv4o+jFWTrp3+Kfi1tfYS8PaejSfr2X
faJOOGXSNf60E48P7ZgbedZAnaII0yTt2mpYXk3hNMY1/qh8aJY6l6VkPnmmsVEIsA2s6D2X30Xj
w5jEe2vHDgujE1CXFJHkCGvCpPAi0m5OAcVYKOUNgvoBIYOIOLPqN1+Ke/yF1ZT38O5ihXfN8eAi
BZaDHitCeDwos0RsbsIcn+TXFHMrjks6uM0L8T6J3F45+rtCTnq4bsdODyV6snwB25IdBSOpSZkg
ppZvCol4s3lA+ZWH26EHtQZJ4/UV89domG1hjX4l4U7tPCboO2B1Ekhl5QGmvPopCs6R8tSgyU7+
ItUvoe/7RLdV/iDoLZu/BkJR5FTopVsdkHUNTa5+nn576GGwNEMgzmbgNW2WzXvZJWahhMFi4hdv
iLHRIs2PyRUQdE+2zxVs0gmvKfZ9J+/ziWs43A/CMDKc8HVu5b69ckxfKcZgtgneshu3D8zPymie
C8jYcV5rlqMAXd9gVjcclQL47llkixgduJrWPuvgxLBuThT7jkKEOHjgMNv4sRMfSl3i3AFvmZRV
P1WK4QWYTszp+xsSKErjFloSljFWO09aBn4QDcURsWR5pE8qcpJ3eT8KXByx4UPeGvHGMWBbuB9q
HPnr8p68R1BcdiGCejhQXcks+lPrm6SS2+ucrNevW8eS+1f6JHkHT7DvQL8z+9tziMjZg/BUSK14
piQ9ui8gBvIRo+BQM9GSiXD5p1NAKHzclqQKTDgb1Pe78vMZUiD2w45DR4arP3bTONzDMa17edne
UwPLj+PGmxqYC+HMw0nXBSAn7AQjzn6TtzdsF1iUlz1lOfr+OCPqCvIZcluU2jVgp9tf97etZrd2
xPO49o+vapJvMjNHtXwpAEvBJBnZ+Mn1HttAbWbmOUK/b8r0vX1KLqfd1oIP71mILm6qoaptJCbm
Re1oIV7RUsJm27A8dg1Nkwx+4SgCyDOruBqZCcLx49OczCGwZDEMtWx6vxNiCAn/CM0aBe6F6hC0
v3CtBTyx3QS5nN0qfpl4Db+PzgYycvB4ePwzQ+3TEKjyxhCAnwcoinR2tin5BOx1JALlBwqAZpr7
kq+0W9sCrVUtDeObnRhspeKkHuYRkzHSjcLrsEYg8p5JjWPh0mRvPZ+fnI8YOoAtgyFgFkyJW+JY
+mh8qrUkEu+JhAnnRkyr/sSobWCl8vq5glAtw/izOhQjrd+S8pc9gEIR8zK+hFFLrcDnB4ghldr+
QRUs+ohOtg5y1qk0oTctd0ShzORaTX2Qs6SAb1aGDVqar1z1rUpMpunp/sjlLI0+54uPUGzzZZRl
/c/cOxNk1yur/3UhQMzBZmsEwv0OlrEUr+JyQXDBM+VxQ+ztImSOnQq75NOlB0dGWRQIgE7Oe+j3
KBfH+Z/c7nOz4SaxYB9dyw3jS6EOD8+qOwlwWUuU5FHzP+aZvm9dWZZko/ynXwwDt5gbTbimJxhe
1RYfwCw85E9QpswJHD4KrVpl/lu1M865UA4GEvA9k05wT7aty4IRX3XoTRukyaYsen1J3aU/tbKJ
oeJILECQ6ALrSy0sNTjrkzHnlYpeHaHXPLnErvl+oKhVsxrYXDCibrNoAdJFv/m0bZlyRDIPzLoC
XAJKY0XVPDlszigDjiG1JSzYU+qtCa91H0uUuqWdywrcZtyL9Ru+iHXsGpCMCVoexn6vhszKOBEt
7xIzv0BSleK9A1mrR8fpM8CLPF+EfR1Xt6R9XkJM3Qt94AT5He0f37/RcWFnzS5ynRBra6wuEXhL
4RaMJowtZyaKq2qDlbMUP41iQJaFNnOXNk6aUAAtZPuDxGy/WFxSIUfHKLG0s0Zm8t28bOnI/kP8
oAg16fqZMZRIIQqx7GKRX63Q4FrJn/fdavYjl5uG2Fd7DMCK9SuTCoBwKUSfLYSxqGR0WfA3NF58
IsBj8b4k4K5jQhjKxJ6AbhpKc6jkF2uFjVZbdpErnlGH/sT1hDRL8bMixPnE3YoKhDPHVg1xCMAr
l628g4tBgxVFTSt7Wq9DfzTviYymgoRe61Aa3zzlMZZJqJPWAt184BqhLiTzplbQIdbJK/NSypjM
ga+CdwX0h33twadvj64GLbP+U/jifd9kT9MuTNJJDWTqnnOyVZS2zPRQewHeWXkfhDhKQ2jTBl1u
2WdWzkqVBbJBAzZJLLDPpfcbD/RCzOD9g15l8GDbhjjTT4yj9h+YG8DiVUinbDvvm6d8o0RAU1UX
u1SWNE+Wyu47BOPFvB/K0ZaKd5Py/3iOujGs9Jzt7eRx41nvB2xaARvryw9EIk+qkuQ5WBYr5ffr
UCepsrpslE+DAUVAPvT8IHkZ593g15TSrI7PPa2MriFAng2S3Eti9Kx9o1RcK3mo06LTfK3liD7e
BgI81b2JGqkbN8a/QCAQDAlV06t4v4V32l4lviyP5cfBIwUkn+xqcVHmPaZB06cSQORSiOg/wDwj
Wpq/IYAU8s9Cn8UdGfpzL4jAaTk+s+W7wOk78OU4YHzNL45XY7cIYmPa8HcU70dgC+KF7qvHXoVa
aoJTZmwUGeBwCRPslGw6ZIMw6QeFjKg1xqXtjTdkmdb8xrRq6hz0Tfutjd+wa6sXdmsFEnK7oyQK
4hQ+U0DtxBwHtSf76yam/zAyYgPr1D6yOsS+ogvIfheLjSMjiGXoE2RJAoSmoxmoPkRiFtf6EFNf
WEOj2tog63GI2yOZ9bDAs3GAFHzREON2ZL6qML8uO2U4SNlCos4MzI71PFpEQIj5JIYu3Yl9z1xp
XRkt9nsMzQEbH17DQHzIPFT/bBZf62l5kwapByay8jYY9PF1cERBFUcMyMlwJFFHQXQjC34rMjIH
z3zJuHgXq33LLu6y82/bEO1hEpF4QfFK3X+WZN+z+3vVnRXTXlVPMz0vmTGs3eyalBqSKxdpnlq0
uJsTVUL0Tc1DFQLgoIrEO8PBTnOM6WPLe8+SgaCOmqQKV9tv/17Jv6oAJNl1HI20DTkJuFowSUzl
Sv45HWm+ji7rPVse0Q606W/9NU5X8QymcZwHMyyYN++ZvB1Qvkny3QtSmKp7FLFxHgzqV05Xx6H2
ooEyckdqTFGXJTJc6xmZ+TDWzASM2PPeGyjhAQSFIg+pp8GkuNasrpGjSK+CW0MYz8lRW53U7QnC
Iu31jWN6t5JhIjsTM/R06pB97INhmgL5kzZVfgzviFhfl/ZmfmBJHgegKB8sEsztZUD34gi3XbjI
aQ9IX5MLvmyjc7d9pHhwU3gJOnH/FiLEibmQ5fb9D0QtrOmEOkoKfMXTpIamIJ2ZOj6Fi3EDrFLP
m/d7ksDoLap6d14+PmYSiu+Cq2m1bjkjPAe1ASFnCA3fuc0SHBbq3xds48UzF7qcBncZz/a+gqkB
qVGNKxLpINXtpke9a64RBgBm/CZgJIyajWMU3FIvlRUtGmTJiGT46phNP+qFYG4iinyyqSsdi+BS
phKNXkcjGQUVfhaf3w2JUqzSUciKyUj/ou9uJG8Y6ffI27xXWEeKyf8zV5E0MgpZzcXI97jJulh/
If6/OnIx8b0XFsyI7Quo+FbVqqeq1DCIc0EzXa7PKRLZVJ8e90RbjLIhKvAxPiYWkzRQDiR5D4jR
513RSnIi/4XsySmAdCEfJzq1sZo4BSILZmU0Sxl7j0G4jOdK8ZY31eOE9GO9Wz/uH3+fP1ciKAQ1
INa2t/ouUPMcocmIjcHfIbZcXBY4GFc5DF+RSOm3JVMeqai9i/ffagd0IJ1eTlknNJh8W1DNHY02
B7BgRfbZMfFkzBT2pTo14s8jDYbyOMaZsqcowcWL848y+u8IF0EDODlpZU1lcvAUvmMlO4khnHTY
CjJgE9iJuD2U77lMxacwmLBt/o6dFyTWrqPkHl5iXMTt0qwF8d4RmduXh6lIYZDNs/3SiJRoEsFQ
jtgljFNRcw5tXZPjafU8XovIWM737ZBij4S/fb4cmNoZCB0zuRo4UqaEO+XXM/FyOjMs2nqiHlmL
7wl8OptddbKEUFZkvrKiPTs2WZhFJK8cXmO/F+CSp85Idd0OcIVbekAy1h2CsR5qLQlmGhFZFhzW
GT4Dj2vSrQm9HX3g/wRs7aUWjRV08ohd04HBTIBK3X63jHzFKN+4Nu5HA0fcnUsuHGERuQWehmOZ
I2AnUDrJ6EN3AniXbZcnYaS4FmUqtleACAzBiHX0SU1O3AyF7S1Om+MTX1fDU+cOI/YGLXXamOOx
TSqYZWXCgVfUTdfo9lY4J9H+1bUqReS0ydva8gTCFNdlkGBNse+Tqcn6olbQJQQ5iHdo5dD17lyi
FQ6KWK6ODApn0sntEvknAH+hnFkOVGYXs5KWhw9j/8oZOpDccD3+fCmfJ9QLlMBKC6JneaeayONb
Uynp7CMzDunNP06dfKnnfO5w6ugomLTmeifjqZdQFSOXPEad2AHb302YM0W3F4vS8uap+sWmDs2c
6jxXpMmc/3SVBG/Phk24qD0STNPIUiKFe3MVnL2RBSYsWxAJnmbjYizh1aP+IbNGOsh7WLJHCMZE
RWtiN5q/1fsaYyY8STBQQ1liwgBYUZfwtTUz3UedgQg6W5AgL26xPJamB4vgYLHt8VjNMB3OqSHy
mswu69u57xVW9GcGoD34sIfdG6gYAh8ZeGxt1k9Ckto9mMqPiT4F/IUYUl+PKF1PywVLi6MWrJPQ
x14m3UPYBRmtoEd+C19b88jLj3BGi2ccFRB20a95aJKVyOH8/E6oEx/2nxR85vec1TnebPBtDBzZ
KFukLQQISJ+Yqd+9euln9lAD8OcrGjk8B/ZK6nGGCedFdrReaWiPuK23yND7XX6Rj44x3bCFUWzH
PWPXmlBuhd9qkyz2clSqiAL3B+fv2/rUuitDAQfTNHGORMGTym3M5hscuHlmkFPloMxZpMQkKLir
7n/Ui72SUJGOxpwMo7/cUSjO622j7kWfbGKErm+QdWK59y+rYfxlQ5JZ2l6cJ/J6KwEo1MwF+CyE
c7VC3dZmV7q8wSmL3Qip8oI1fHbrcXX9Je/W1Ex8CA9/9X1AriK3QlGbjbGbt/3UeXSKjKXVSpf4
z5p76Dv2/4BE8dOdXJUohd0mZJhHrxzzExPXKjgU8viWJphFzxPYUL/fDVOp9cr0yMqcb/6fq6HL
iqR1p70bnqI8aGD0iSJjnXx3t+14COpSuiQOcwPJm2cOmRWAxSLf7LuwrZOxVALKWNrwx0EEanjU
j41FvCDzzM06ioHzbcKQ5Cub7VJ8dab/RmDtDNvo48jOplbCvmYYjQ8Svv3yWHy2u2LxHZqtbDlo
wmEqCSuXO1Y7rYE1Mx9M2FHxpXs41aWl7NdWplAeyr5XN0xvm1CbSSSN9OzGgTji4zMl2J5M3cT5
MD8Y3QVnN2byFTcnYPB6LlN5Xl9x0vjBe0y3NtXJ9qjpY7wkrh1YrJQCeH/MkqoV45rWIMW0xQ9W
DkQvsoX/U0uR/komGznEjW60QF3Ali7UKmTCTkeEc5dUY4xNT+0Bz3bFjd47AXrBLWvsqXwqWogD
Q5uL4J0gc1nU+fYSFhLaaqWPaTgnXf3h4Ojo56LH9/zgv1KlSzQLrF5sk9JTNERzs7PhtOuExhax
n4LMqMzp1ix/riHMKakcmTqRfF3rP7bui8tu9n1wsotDhCV2KSEi73DsmBupeOKeNWmrbTXOz+1o
zemKBeVGOx10ZcISytI6eGHo0KkdvOLIq03XCCmZAOb6PJaCX8t6Q/DVK06w3RDFNCBEi3m9NXCk
Hb11sxzXIwrZdPECaO+oGvk6/bXO9N4nYrkFW4h/0lDK1/UOVrGJuZOr77sBfWhAEji00202VuHG
hsRqINTFYEeSYKVoY8VxcfvUmJ9uE1t/awgFpIda36NMUawZ6HCnL+X/PD+zkV3gvFNuS9TSa+0x
o2XEy4bZZDgKuPSv6qhNWF2p0AAWYL3kJsbeFZTNw3qWG6JP9+iFPw+3xDO/Mg1XeBTVkfpFFmU4
jK1/3x37Fn3Cu8mV7QX1vN8qaWWHBacOGMJ/TDZU6qiN8UF5yd5R+VJ1AbBzcN/O9ofZ3YWPN+Qe
+X0bU9qFrzKxbEaXgH5uKp4etr1JQ8nfBSLuQJAHoZqsmg2bSl31LjYtZ5rFjrNQqvHb3M6UKiT8
s9WtsJvlSLybjxLWTtInfoXncUKVTGm97jWgBEGYWt7LDBsNixQX9BiZgxYzCLQhoZuD0WoZ2ebW
fh6eJ6GByK4ruu3hH00XrDEGDnsnfjIdpXrrQ8NHLh8NNKYztORsXya+E3hVRG3xKeWu/3cXmlBw
zcSzWCUZxVjACh2h19DURG0aaZPqqqaNvYwnqHF/td8RuncYbyI8uMOI9y2iSVoYFqo7s0agxwkE
40VpqAKjVmLF93YU/31crTqwD5PIg94qi9xCbde1Jn77YHVjOcpmN5UHUyQufMMA98x5E5ugzyDl
D1mmlQfbCWqquyDVvDslDEAT1xfZXChSMUwdtIU5TueFbQs+E0ZU3i+hYz/Ys4Gmz6V1qFi2CTrb
PMFpJgMoW3xO1arWPHUqOo1p20jroYu79FfttS9f2VD+9M/trbmc+78CcgZlZh65yyv2RajZcOAg
5f4AoQtbdOe7VWh5lRjKqvtJ8OjZ18MqKrpBaQry7veOMVY96CHr4JyK3TY90tXXiA1v9JBedkhT
MM1PTHo8Cj9QGcFeXuuiYnSVR+SELEZwkfZyF5XqWczQ5+BPgw+f4rRTRhhXGyeXdh+saRpKGrTI
ZzOJ4lQfNUcac1Iow48kKWEERuZRh0sAsqoGRtg0c9N4whLX3ghR/fi1nqrW0H+RoD01lbQmn2vW
SiZgOwA1ONG1A0juTIXSFTiFEKCN4Snmg94QuMYluzHeW21kY5duKihDjn/LMSjTDTWkw0Utrqtx
QEfSKc4mIEp+XKbFgyhMGs7FKT7Lx9OCMUUwdoQ0IYDh6DxJ+uNwSdYwXoP9i7tAaPt4xwZR9k+B
9mMlD5dYOTpzUM6HM3pCQD/yfXcC1ukrWQguuNIVV4IO+Id92E/SQugRRZvlAyZ8TaoSBHkBCWQ/
0b+ZBCtaZWFpXwImW8TYRmDogl39b/cbkMMzJVy6nMvzGKI+kKySc/ngzq672bzvt8py448ul6uh
NLrWA9yCJkQV3Uuulfv4vTu+4HDyqiT5fcdLuWdr/p+7zcnrkaxfFPRxaVTnM1fj2sv3lWDwEiXQ
59xHVguXzLJrmr2Kdp8rqMABrjzu9HCXpzBS8/Sv4ghy7whrhzi8BJbtk3xBKks906ZQPE5ilFTU
zZm6gdiJQRrGJTEpPLBG5sRD3xMksgvw/eM/s30kBmbant6kllv+XePhnX8fiovwPIxRMcVYSf+o
bSrQXdvwlYm6qqMdSZXEZeWSUn3x+9p+9fbWTsret3cBCQDfCqhpl/i06j8wBCoUif55n7wDN8RB
AxYo+x9Z2UPP/eTpXKOnyUmBVNJSuW7KPKBsNofRjzf42DDUrALxyVduZpk5urJxZjSJgNqoRs3a
wUkblkGeiOqt/qSBptCE+RaN7p4/09h6twJZLGsBd2YXPdSQqPCWJ3ntvth6xsRGiIL1c1/ViCs2
SJ+dftozbWaGAqniUTI6DEOCqp2NLSRVoMWxw5rc1hnVkUmck6tk9gtjlgFWRFnaFDPoXBtAIN/q
vTwpB9kS5PoL1pVVNq5RC98pAnp13/55EtabITq7JSJDBM2YzgG26eRIAOzxrwTWHlGaW6GvatB3
y3YaqUKi5CxiakRBh8FJE9HKodJuAWmp7WMaRmsa2sdWefVlqxdrxkug2AGmsefanQ8guooYbTKo
eDJ69ZrQsIANahz+Ek2UunjtO/WRQoDwRy7MkBWVaH+xNWPB2KvaqxuINuLdQ5Otbg/gWZaihSD8
TUji9osIiE9bcV562njElWepvlaFQv+E0YHwyWt5a+GW3dcZbJlSAm37h4FFxBcn7SQEIBDzJXr+
MxjYt56Ci+98b8w1dVx5hVHhm5PB1kaFoBIq4JhnkLmRL9uztpZklzGnDhC8z4efcqax2Vylv6On
mbWtmimTWXJn8RqLxGx/60YJZZHOwTwenw4haIwvXhQ+zX8Af1tK/vIItiq7UUpCDZwWJ7vNliBC
Oe4ar8pwijR5t76iZ7oV2VMc3PpZUzFqFd9ZVNTAtdwBwhz4zGd17I3cpAVJIkVkNG+yeUVdyMGV
twgMIYHMji7tQopTFdd4zUrlbhWe5Lhfts1RUMlLlPsb91X1RMrhuHiF6PFvQyYGMY6aZCzL9mXG
mDLEyWrn0R+73pZAFS8YlV6C4H2kjZFiQsfo98RMpAEFZxa7uhwkgnRpflwZREJEcphqf+XvEnub
QLIx3E+pQiXmrRuJZCAlM7WHIRVXr1lTxfY6SHTSyBfX7JpCXt+PuYbZu0IeETi35TlqGs+6wvu4
SX3AF24oxJGGi7LldPaJQz7T8VLAHgRNcv9xwjyb6FubHjitOxI8d8gMlj6U78brzAhPPSlyzFgj
AtuLdzYpaibiTE9GabjkDAnJc9FyOyGqT1fPE7BaH+mEeZYTUKGDJfHkvYwYKJ8lJwQV/SThCQ6o
3piW7WaOFHC8w/igRMWk7EOmkzOu3r1r1dJldY80yms/OXt0w8MzgxwiRTi0ZDAFxlA6OsZ7dv6z
dSsX5sK3oy5Fx2Mipgma7wE2dR9WDPZ95yK1le1r5jIVBDP9MbzapGMKVMvdm3PUn7i9zpeMHCdC
8Jc+JSASZJEtapc4e6M9BZSHuE0+1jPDQdazosXP4DcryZr54G3ZoRWrziXCHyV/RSjO17c2uHyG
49QUA2BzI1tuiip59vOsukaIP1EQ8AgGTFp6408XaLBk3Uj7/L9kQFiv0X1jTWsUfgvakzQ8x6QG
3zxGrG3cQa39zYBn9SJMOuB0aKexozcDOXfq6+1s58BUvoXeBJNq6qgtV7ynnDZy8g2x49iqq6pB
WrIZrVHdXJYcTWXop44adPd4l0kNUcjAtKK7jTa0MA4naYeqLg9NlnYGEE3RqfdjlXsRozaTxxtm
931YgDEaWWm+xW0PV+tjVvbEdxdCEhvjJXktKHL7d/QTPoebV2aO5/YPEY6Ps82hZY56/CESOKhP
2O9gRHM0dqopzi8e+OF8t4AD6Rh1KekIvOQxpkegxWIZP2RNUcVAXJLe9faZ91t2PU3pgUXAFM0J
fk21sOmApxk6N+d+3pClisWyvdvBqnz/8PQVcjox4uJMCltteF0YsUHddSECgWtQXEGM1eR7bbGS
Q7UqfZ5qq1oejdTH13nBbT91a7BovL7qHcskm+yUJsFTI89VUilE8Jk0l7v4XH/kUn8t9iOQSO8x
Q5+Dj/vtI3khdSrIHyeZORir7gCHmWNU1z/D56SVeFPoHMNOqO6nm6lbwXDsIayppTTaxgftL/M0
AvNqptWeJoFVEaX8+IzLwqqiOBtHEpap0KuflYpOwDhEipn7g/qLo4zAOysQV3B6EKZ7rDYwWTSr
PELCUjuo/pPWMWJ1e55LISZgJCTvyYiQKzctfnjWT+wUrqJyKYtPSbQ2sjXyPJbi9lUKCTpKnldM
JUpNxlKL0Nor5pr6FQzPB8Y8B6s/odfV+DkTeB/SC03+oHvz5fgmMb6BUv2l877cZb4rSlbm+bzM
5lsZGQrj132XMEIZumvzJhrtUsxD4azEu2FKT6MieFaDubXgtnasvGZBCGuFP9ys9J91alDc9W4z
p5RIDHuItTFi0PkKkf+XWa/a+dW1uttc6aJlnlEdOY12wPFaDD0VXM4tL86YWiZk24dPZsH2N4W/
2QlDoshBgwCrugAVL9bUNyVW7N98vTfrDv6VQAtMS/AEOw6IbI8AWiabaYGmTaEMyJNiJaN18LQb
ZMYY9LFxUYCYtuDq2bqDQobnzBTgZo2cyKtvy435HIk9+yUR/LtkYqkmKpUTZUOef9RyWWv2UpsW
kV4N0zlqpwfqRZTmEeFwICgJ+i8tBfKAbi5qAxg8DFYGRbn4/x8IJw4DFdQCGJaRlteblyAuAisq
mI9hgzUOO284GJQEpPeWY7D/WoA4A7iDuh1Er8q+HcwpqfUKRThH1GEXH8YwOzn66iGp/Sc5J9/l
360vO57E148U9u9aX79QTyrbFDQVjHz+1XrfyU8yaQUA7C1k23NxtvnFaNxEN4ZTMcJpwsdtJ3M2
dvd+k6jvEVuhfoOMfgLEkCV+wiawOOpfXPKDP4V7kOiYK89cGjWH/Eqh22IkEVsLK0+KKtW7LpK0
GpYTikD2btbFlWTljHdrrfYwjaIpYEnqiYL/xDGRQdmXh0YBK0t31nHw4hMGk8Ojrv19RrlxUol0
BTL5SXUb4RtLbPT0guqTiWoIq1T63twSIc8keYqiN4RTvJx2PwG3QFvbUjkp3wPpXojKLFVnE58/
IlcyTv0TPKlT0A0ZAMk16pIg3Tz23/adDyQpeXGp96whZnQW7mNIzWWTu+I5Vr2M32AoI2oHA0Af
HTIZoqpI2zZrY7lCkQH9I5V5qCdydmQ/OZRiz5G/S+wmR9SDa4vVK6bxUCWswR43tdoAZ8nzCRtA
Ko2OQLWCrqZmk61HaMyghu+iihgqXm+68H/ChGHUGtF4Avt0ZTLyoPb0VxaOKb0YmynjD4HqQ30+
g0/2+OOXyxO0CGkxWgm7Zw1oeh0JvBqJSz4z/9isKMqRoxGDTbq4nyy9NrmPtUPkPTVT3PcFNHae
7uhrQIUn4A9UOLmvVwGc6KmWu7h4S1CjenQPR3Orw1/FHgg+VS9wZ+LoHUrLGBBbv64gBsSsNdFn
SnPg2IABC16H6NKWAPKNVJYhUccZ3nbnjhy7KoMB4rHuhazh+/BsqLl7g5qpfndEziGKeyfJVYv3
ZSGjCZTtwcLK3gVaVPIEHGWIQ3dmPqGc8KhGgWfbsd6ubnj9Kx4DQzCemqgBF1fpVc+Bnhr2Bkrg
QiOyd8+fjAACxPGjnyb4TtuqJwrTwBBJJGTZtku6DaMbig7IwDQxVZkO2Xm/vwnHCaWM0FTB1/xb
XuaRUWUk+0Un2BrB1WGbMxGIlbZIr3wyqjU0fAFUm0ip+wRSApLfVeXyikBDz7v6VYaZo5fDUbJ2
nrim30kj+s7tOohDlreMI7upqKbAKknSRXWufwdWdTTvZ8WTLoGG/++TVekofOGBSlTnjZAFIz0i
Y0VUuImDUpkji9Htgl3wPO2ScJra6TS3PPhT7nuEMeb0Pku7xiEOfc7laB/pbTP3RDb3kRkB5pjr
qltpy86zcC/RS0jzMnGZ9nk/BGZb08d/vcnsXe8hPTJFIT1DgpfGbTX7eMpI2Dr0JAVzFK1xSU3z
0AcvIVtrydmjuAkZawU8ECg/9HPCVVrbtdvivobp1tJNCma6r8M+41PQM33Fy+bTbDnMto6Db764
G8FxnXyo0dYmE+/WOwv0XRdEwibWdXDkES1tdXin+KL5Klfq1+l6QG0aGGvcHYo2Cpe3LZOclmY1
ZclEXlxFo32ps8jtc2OOqe/xQWJbRJdixgEwgNeOhScxhynBXjOdfy/i4jr/8TIeg+2kMdZ7tHsR
Fkk71Ky3MXaAVCJu7Vr6TQGZdpDiJv90DjE9GOfLhLTkw4YiiGDwJ10navg5GZbJi0+qIR5ppkH4
ZImUB9DPJlSauQFBMv1MpobNm37m2VjE1oR/gPjmHyOTPq5FdgFic+6oV8dUBz5xXPY9zaJp5lb0
KI7XYwwzP0VR2NFBu24syTZPyaV0TflTMHuAr2TePgFh+U/K5vmS8AtmxOVHeTJOQm75peNXANhp
zRqLs5LBu61ws93DffpUsNPIXyrF8ceOji8m15//QkTmj9dUs9aWgGzDjf0q+GLoeMLv9kIIe2iA
A6rtggD3v6T15jzU+/JuxtNK7q+7kBnF8PmRHfmugOrd7dbRxA8WAuY9PM334F0SHk1Y9uXzc757
XmjxSgvERsrCXlNkNjSnUJnHGxUaG6nTerjfpcPd9dfMQi9Q4YwlHPC+wmKo+y1Rvt5YsRxuHMD7
CPpj1e7Mqdgm4UB+vguN7KUihjAuZKBoojm2dTmOtCYTuR80/p9EsEUu2+sQyQtxU7bHY0bQ2NBx
Gs5OvqwInyZkW10hVr8wxevtOwoY05uE2Oo3iWNvT0aiVIkFRLUvJgrWwJ76BiMyAWPKfqgE/mml
a2cgtrwKf94YSsHn5psbkc6pahvi5D3GDEezzBeyct0c6hynU4RW33m8wU331OjcLliNaKozipDf
eAjbFg2EczUgcF/Od/oQtfrU5bEMJ4qlSi2VJIBz6K2oUD/cR8KT5ILX0BJT00Ou3h0Kmcgx8Hee
7bPPFbY6MxImLaUh8upDUYJ9jMwtjeOoMF8azlHJ9+vlU/0I/5Kl+K6xNyHB9oLOXB635OCUNPVH
+aZU0hULdbdgzI7N8wK66AHvFAC5HuvNzyZhBjN/LGMRv0dBfW77Os1jZd2LQD+LP6ZShtT8tEs7
zOz30qgMWteNgw4Haz/r9CSsXKnTssCsMVaHFKGYIAo4wge7fYAgkskobAdiahV+QANRWrJholDI
hZosHsm+tAvv7soJNjqFUWvnH3/6leam91C7tfWWKfjWdVQOybzgXN2pKPxzkwTn39gQ9J7CtJ2E
v/B7lhez5t4IG/KSlDiGGL/3OosXkty2n81y4cuuL+PpKSWZaCpm8M0SHKJZjeT7KJ7dBHy+eAZ8
jjiJ+jhr6PNPa53FCP73FRpTZq8sWGseID7iDpUsRyysMcPyeCVzX2tXO/I+sYcIGoy+/7fTb7X3
UPZH4Wry1ZL8UyGgJDHQPBxQfrHdi5a0NAG1OuGnZF8Cn19tZIvXrZgL9Wa4SIoBeL/5wPxENrVo
0QP/rVOT6vYNuEorFEh9GwxEBHtRsylaXBSTd38Cz1lWYiEhXkWO8tkdwJ5DnTJM10s4t1sTGKUG
ad+QzwC2+xQtWQI/NOxZrBQEfBe1fS7uiT2CzrqQC8Q6L+dyRHs5nZQC+dLMqnkbpT1UXjeM3xli
zOGjAtFA5dWnHphBMkaL74x1mmP09d6s577mWf+2hGH7TJ3rdDClimOqABv2gxvgJN6Be6LF7ykK
5IcVrjIisBx3fVz4Rr7/4Xd2o0zHiTRuGLwZ6ZiQk5I/6OIiHWy1PNFQ8J3VsEoMcK4GsgQnvHao
5qPCzubt0VuM7XHqYnh1og8U38wWjJGPxyJ0c8z3dQKaQMV3Ivoy+U4QzD9MNWnAgjuVt4sJntX+
mjIcRCydpeI60VC8txQwSjjjZB9WomcdCb0i3H/whkL/iAOaUOdW+aska0fDhs1/P/5pwNyOIHbj
ucMpVJKJ5jBtdwB04ETnmgoxBZlJq8895XnfTTGWE6gtuj05NUun2Di0bbDnXBsfUvaGaqyS2EL4
2hkpGaMAT7RMjGe35h0bR8xAPz/xaOH1Q0mSdjyIQ1pSgATGLcwvOKFpD7jEOLwjMLrvQ1iyfsjk
wWuJwFiRjNyDD9lx1wisyfif1fmgFvKZgxc1sl4x33NaOyq5cL5VZJ7x7A9xx2Zmpc0SfpAkkPo8
fv+3kNueTrb6wpgE3EloVDjP4/A/v/OgGoP/E4dedYR3y7VHDi+hU+234li+9Ni3x0CZvS87ZPQG
nOOhdteQjWPot/B7vjhZLdDUnAO2ZqEeJvQLcYGegxd1LFQpb5p3y9PBwXDgQbfeYvXkq/TFZ6CE
ti1HNymIimjXYQbzMNZcBfn6RCirjHfhK3+R0gZ6GYEDqGhMC1pIaH4QXe79nCzZWJsKcF1AWJnj
VVSUTdfdiKzhpz+NkxOo8AVX0YpUvYQkrJOXwVDI+x1V+bDrMcoDad3QjbZ8WaTzEWL0Q9c/Mjuk
kSabynjsNSJiURsZ4j5w/GuPiDdtC33Sur5sR2Ho+GjwhMQfWXVeg36XNbCukYXuyzrDZiE6HuHe
qK00bX7s21U1FrIVNvoJ4xapIJwnbflAAgfBmBwFPm1CMruM4glieYiGPRiW+9Q11Oke8nQRSqCw
8dtMCEtDnOsQUPdvnC7+KFopowXFX4g75E8C39W1k09CvhXRLC+QSUlUCzvqgvmVKpS3w5h8/SaI
j9jMcCZdkPvVloEEUmnAsSfH0T5rBIp023jeK2V5kTZn5d+Tb+wPz5JeNhKEsIt7blQtGkdcYUWt
Toz2RlPcBr5gynClAAeaID3pqm7mvmDaLT6MYV0rcdOd+5oijc4XS77Q4Po5xglrLWHC4snwUmoi
GHqOfvPYK2kOyrhAo9RdovwYaxTCVEXQr2NyUi+k/pL4ivFdij0sB90Y6Ow9yP95JqEI/NOgoO/K
1sPOR4GMjilCyuLZ20M5EeDlvD74wwvLZAf9gVwkiZTWM5tsaNDVvIAJNFLarySOKbXqAK/H0xao
v5/x7VjxM2cEo8kjujkVxgqIm9CmiPj6eD20A72opo5xFw0Vx8UFu599JhHtQKk1yv3JPYgmrHY2
nHJ8KTAUzNSVhm2PPaS+fugH/F8oP39pJWD1AqG9kNAccOaZUc2Cn13mmM6vJgcIqMLKPn+06Ik3
f1GS3wUkNmYxiZYCDeeovUXx9hKz6Axdv8dBIGOImToXY8k80SRMCR/VYrocWR+TnR3qtBWMuMLp
D5jpzEuv80SnQwEiraRjedKGAZX3jjMSdpSeabv3dGEHguut+eEDbYL4yH9p6nDMHbS+2q+8VO5Y
wioHoNONDV4zkkTfPTCESlLqeeLw7PaEPy+v7Tt2HaK9QeWMFi6MycUDGzl9PGlz5t2d6MKVMjio
0PsaVGfuv1cz3y9zUxEIC9E9O5G1Q3Mu9Lm9oikV0GyY6eL77mJ+7S+N3Vosrzohby5LJhFjwq4G
H5s2bEQybzOlE2Hxz0giXEt0Tu+c97nuEXD/Hzin5gxUeTrIEUQ5slm6KYYi/buaiXLSUMvLz/wi
RGvSGsbrXSh+I/Y9HqzO89NUhJGBZ78O5PhvKuO+H1GIoY6lUbEHvqNP+HGcDOAlOVQMOhimIWel
n2LxvNxd986p59/eqF4Z0+XWEDo9Rsr9mTLRvvK8pGJQjg2+rh79MAzDoM/7mzjxIV+iu7DkaZ7T
zvQ4zIsgn2MINEFdXzCuE3ZqoyryMM8TGQ2xvlytFLbll2qg6NGLkOPuOZ5Hk1r6KGsZTKTwr3AC
dlqqCxdULdHjuxmqpX4nwgg4khjwj0Je+czolKB83TZb5Dif9L3NU+IbafrD9VvKn3QQ367aXBv2
vZPUkxirPzv3z75K2RbFw8VgIZTQVfYUdCn0mDo65/8s7PLAkHGAG+vVqI4djI5PchLRmEPjjHTI
VXR2mVoRfWe0KmIWXnRiMXIuJM5bVFkoMoK8j8mp9+CaqUmW6VgfG10UiG9CNw83pyByh5inZxeW
BH1DfIsubsTL6HKa2Oyd+BqwcWnIj7gJbX+6TQzUYVw0HU+QbO2RKL914GX6fBA6hNga9TJtTWrt
ZqveX+uq/IQRaDJKtBwhcGReQzL/RaJkRqGDaMZL5YVLueR4cCJOLhoNCMHmSdcQG1FX4bNa8D56
n+gbeYUvTdIOJPR0IROS1sf3H7D5sdflCzqRsB/QmfMSEx1qNTaxkYiyAuCTjH8saxhgH4rKYPmU
hvbv4yxdy+l2Z93NHGQsRMAftw/W1T/y4TIG4T4dnmF/cGS8aAE9bwh5KPBlF1AB3yTFarSZhWep
J0EO/2aoKDa1YT40esKDOrGqIqGJRbZxbZVjEbq7/S9yswHnzxJhr3NxZk61a6zgEidLVM+faiZ5
0UKDGI1qvJRqOzqEW4kXGZgJBU8SLJY2bx5OntSFYxcQf3UXIyTUttFMYMYO6sPzF1Tm8tPX+Oo6
a3eOQ2FJu9qaroAd3eCDBz4WDJAuzIHFoAnD9nCZXHc4IFoAPafsuvhQ1/egxDaU9UpmJ5nwIWhX
PnsLnKK0zHlVtXUbgPiCe9c0YDQPLgKL/ais11b0EckyPJKirQ8+j2BC3OX1L/4tyjfD8lOCw+n+
dvSBSJ/zPQNm9fDgrnVRNLI/iPXrx3o/HHDSrE3t1CURbR07305lGJh26gl1qi8/0xSkZDlxVxHX
FmbEqjzVmD+TW3DjKNfMnvXZMl+1JC1lv5lxj3mrB7rHPpJDBkSiC89JSPo6MR9BkXIGqrDtxZ+d
7J11thh5ZES91pxSe3auyo9UWL0eIm2SPy0nWe/XEG9swm4x4q9WkfhSRNbDeEGqj4gfBptghHV2
K4/5ILLVS70iIWmrggZr27DdmidcJBajhLFNdo0BaPPRkQEp1jNV5tlXMeciukRyLZOx9/G0TcgH
xoyvaRskBpWkR6i2y0Oh5mtnc0Fh7+KS6qIAD4KqeXq2EYIwbiFeyveZ6xkLUrwu7m9EFiM+88gV
mITiWxFkOGrYHTdc9TduR3HBQOKmqm5Z4IDpmhNuKtVXbNPVrdTTx1BWOdpngm7hq4s3YvzNfjgI
dVNWCUORcdcwNbqo2xz580JR+3JiwoKeiOnSIrDiqWSaLVT5NYC3ub/t0KBWR5fKq4AIUcMunyQS
30B6U6hfHHKWpac61CLCgZTIaMxSeJhz7/SLfibBomcFYRHbEjlD0/cE+uibq4LbDxcr/tRAoJrr
Y8wVdbYI+Ma8x0FYig3WO/OP8q1CVPS4UtJkV9R2Cb1L5VgESnNxna/HTrqf1MsMzuxd2XIZbu8E
7XfaVjVNGi0vxR/ZxJoG5OxLLv8mtPonux1IVXY/6J/9KmVZi/uDBl698cSuNhuzpYGXjdjSOJ8W
2ZaTSD4ZmwHeoXS6v3XFku/tO6ebnI/hs07KlrOmfBy+2um80X++C1QU63lpaxS0Oy3xV1xTha1G
pWu6hnWACpRTq+lksSMjV8dL8vAIKhl0PRKZLmp+DzF0bM3Ljyn+uj+wqPo6Px4qRss8GpC2fMLk
PXh63TrSKUSJMQmbe02IIAHy5a2pAPTMf+DIylvxGBsjgCoUZ7O0/t/kwXtZihesph1e3BDT21VH
CKTL7JJMM0v7fauFeARglZBR4vEMQUL1+MqfUQA1nAtrcgFRNElli/58n93nR2e0RtSn3gZFekCJ
0uB3FEds2kTgIghdPxDpn/2a3kcuOt/f4ijPb6u8pFGVKhp8yN+6hldlhfOP3eVyx/GKMZxmsAg1
ZCTAENKVkafkgk3xPxz6KeffVopp4MZPtVPm4KTp90whO+6aTvVbnOzDZWpjBnGZOiI6/HUkMMCQ
SldLYmtSNSkX4gYcvXC5HWCs1aebzajnTBpX3C36kouJznMwkXC4qYXY578jA99DDK/vJzgijZS0
mo8sg6hKrav0z2u1AmyLXd9dBxohmdhGtuWj3cnDKBj75lATorJU0zYBvkXgOIrM7TggtFjose0l
Z91Mj/P999zybX80t5XB17UVMNC23YsVwxj7lhatW8bjA4jsoALtj0VlRBAH+/Hpe/RJVf0GAY8+
JTPZ+GFOBoukSdCO8p24mCaVQab/m3ImoiS6IFudDP1r4WRTOTV6WBREgGEzUgiS4XpJq7Dj2Ci8
Wg+hJKQz3/P4hB6iv0SR6J7n391SQEcDFZKOAKSOkbuLlaEg9RbG0nWwtoU4lmoROe9OwVlEMmEr
3jR4tb03aUT2gRcIeWCf6BSy/l0T822uZdzx5NJvB9erPA7Y5r7ffgmjIvWCPK8mPaS1hOJDWAbN
CXTu0/3ul2vZdogYx/U+dzb2ylqiZvqdHDrns665pokcdphZL2vCgndOsNHJD6m5btR61FcN0bER
OUA8T3fE/aFaXiw0Z8Q9qziYxByzOpAW4xRXBcuKjypTbptZ3K/c6YI9LMUDJw868zgoPytH665t
exxSu9TMhUfTi6TUp8Cjc2X6ljr14cOU/n9yv2GYejJ0akmvw4wQID8XiDxRYmlDtfCLNNZUB0s0
IeQx94VIAAcZaDSpGcTFFWQs50iubB5XuLip+l6KfTW/sI5y403Lr4w7ysFhE5h59YtMO4xSMpg9
hokTEs5XOmanpJHFfrz8mrWoyoaG25QSZ+MU3/eATCEovh8YG1cZ9zNPzDf6BGMRlBexdu7Kci1i
Ml7V6r22EA96tBL3L4of4QZw+upEQ4gss81lRHWD8XTNZiggByvKZXxkPndCQ8m+IiwUGmGTgJEZ
BMO6v8/tvTYScRJppPYagLg3xcLLRMYhp39a9cP625Xk/yCws2CPPcqc9ldL5fsdnhKtYsHRYkMg
Nh8RlzLX9k0X3hmu9QKPlYG5CFEDymo67Fy/L9YeStIJXCvAt/B3vK7MpqtMoDPaHO08j1sKHg6s
KW8wJ2z/Azarl+RED+tZuY2mAfXU0tJSR0UVfqrdrSIpCaBb/R1+/ulxsnxgJ/pC7TdkSxPVKKKC
QtdTig67Ns2Z+1Qz3JPFC+EpcLPlcsWAdnRa4DjX6yNn0KaIObMXYDLS0XuZ27pHRX551U4FeSkr
PH9AcJQ5U/tmy1dr5KuymG4XgNAEipqbNKZ0+PaIMQCTBCVUm1QoFAnS6Pw9KC0qPg/d2OSmLElV
BVyMyOVOsV/oQOC70w1GfKzowr56sq9OAVjveZGKZ4F1jzOwhCxTdBe+cpd/AdIfPyKZbZ059yDG
xR5wJwDeWNDNy6QYWDUPfvesXIbX7G/aeKzZE8ydftrkUFQL3ablEvESlTx1SnJZDkCsM4e6VTaT
4lTjJBW9kmX9AEfqnh7IKX14WG5S8+oqEPu/TGt8g4BXDjigKOV8CBJm9TiF+LAm8AkqDDSQN4N4
N9mlY3pWVp1WWvE21I5/ZRUlrVCpmLIN5kJ44fx2fmNkLTcZRVq1RDPz4+yZC/BlGi5zrC577YcN
wrJGLWLIm3hgBp1ANbcvpj9G5yzH7GZD4WbfBcPPtQmkY6bVtmDOLCtAltsKv9UwlWKFhUFJKpb5
mTfCtYOSCfHfWSjOU8hLrEAiKiNeHeV4J/nODL1h9fZNtDN5npWBKGeIWEFS60Yk/x5t40FYkXbK
NG1LhjIkFViglL2h0c2gAjhC39ndFi/MXgMOpLO2Ed3fyAgNogOqv6P09CiJxgNry0U/ynxyn41k
VNdWovQRrQ9GmOVY3FxwJN9Zx18oirv4XgaJjnPnqP4QExPId4bKe0UXHgjQ3G1B0oe3JvUIllL0
OBjvZbp9u/76O8XKtRCi/KNQfyAU2n7YkAYqB4zDE3Tks9lMnuVglwpR7esg7McKlpTRN3U0+Mbg
RXZhG4ZGFEYfU7xNLCueSH+4YenCSg65ECDhocFAAxMZFjHKRU9n8OeVg92LO+IWhK2MUTH0WI6x
ya++Xibi1x+XWs0V5Oef4BaEAd5X0h27Aq1YqFN/SAAkKna3V2+VS1y6qMOpTiNmJy9OEIOq2uRM
GrtTFiTGzDr13EXE5tc/rCLF12YS+00BZK+q2Aa/eKcKAXDOsN7QsqCmvC9Ze9PKKC3HJ1QJngre
rTb5XEm9yPaU0jEQavThZz4ZZ1gvJUFODwo7XKkx72pdZBhKaM831jW3Brl5uXgssCqkhAwARZbk
kJ+4HaJTot3XIcGIWe2JQDNahun+DCPgYmrU1YtmanPJtaZCLQTsCjmuT/efqjJJKupGtn41o3Xp
xjshnTwaepCcMVTjz5/6F2mEJdk2hA8qL3sEL47NqHwltDndQFrw7d3bgpPqhLRRZAhXSPiaRK+Z
oEM18k/RW9vUWuxj0VDjuDp3+Fqu84sgwrlqq2sH4qZGK/L20UcTisz/SWxQInIbfqiaWXr1sBg/
ZR1YIASiWuMRRWRUeiMepnxA06uuFPS7j3r7py8MH92q2LTmZ/ARbZ1Bu/l4+ZfWLoHXjkScVg+f
AHdEBBO2DBG2MMBw88oc6TGErdrvUssGGnSRHJFoqka5BZ/+ubVGc6R+9n248Egn6Z/mULEV8/L0
WBe8Hg8PKlBvXchR/TvrpGMq/qqaUVJRVLQU1n681FB8EqLRZas+zi9CiDbEjokJD0s04+sSRAJw
cbwLZ0JvreP+7fjzTpiijgAxEsrizdcNlNkVv+HZXtlQY+L5HO5O7Jtvgpi/LWc2lkdEuLZHcG1a
hOc6U1xIqcL4ZLbObJjf4QbvXPPgO7rZvx4ln2eeosNLcAyadaFIjR/K2Lam2j/H/u7HG3M+0xg9
NwKg9zpWcqGoFiLBO35d6jn32QOaBCkfFbDljR/dyTHxaO0lSyEQsWet+qNd2IsRSVurGpmchM9V
uzy+a64wCEF+R5WP8uIfBNwcabgO1esw+4A3KA4WA3CtNuISHgkI3uEdbru37SrFNvfRTGRMXHTE
D3L3M+DVLiNLUqRY+b7U8NAfEm4Uk2roX4x57R3hhGfvgvUltQGbEvcsa57DuCMZOHLtLBm7k61R
GJR+UqZW17feEsMXZ3GQQGZZD2XAJ7ulMMXNmBxzgDJMFBL8u4ncRr0MsXjdpXiiU0BMS9YExCSW
atXigX8cYtYX02dvgkPCLS3ZXn1Xlpdjjkw8AvdG+BZhk6JffWSmWIwHB8sQaOIdhxY0JkULOm4A
qMCeGwT0Ub+/QvJNy1up/yVo2N5LsgbK3uMMSooFwaGvUhaOKAWmqfRVDvejLgovcURIhdrAqnhE
igdqG+rCwJl3+zEhqWaCPsYV7Wt9r59RbS+ddKmsZ96Nf2AuEckN/Nnzak8y8VIi6yzHn0IIenCc
xXQCqVy9RnZvc6odTfOR3KqruOoCvpQnjZNGq4tTf1aQR8Ew+4pHjCWQwIkCYtTSy2X7AXL1Iou0
JUFZxMOitbHU0K2yEjZ28bhaXJS4bABW22bASU4daYz4Gg4Kc9BGyw7CICC7xW6G9VpWi8QhbimW
xljhAj3hggAndD58TQHAFm9aVoFbMA2Kt9ACKeS+aQnJaqiLuiS4+jTz/vFbtHQuO8+pU30/VjKf
h6uj8ovTREqeIUvVyI8EEKZ/8aNh5braYgkoAFKsBVbeC7oCjHIz4XXp8s89BcK0Ci0zt+S1Nmuy
Wz/5Kh7s4VQzEIPsdFgBK6Gxu2C60rGNg1uW/Lefp8FW0K+/FFXqLiFyLGjJx4478VwWnrS+N1Er
sZOUDln01GTMcahD3U80XwmVF8ZM71wIs7mpCdIEe7Ekn9SizHeZYph9DNi4TauKALEcY6AomgcT
5ufbOX1KtZrlmq0TblFTpQ47OH9RY7Afg+ajIIpv1R91BKVrKJ7KkRXAILKA7X9mLD0Qzw7tHh+0
IugOOTe5q+JvcPSfTFd3RllSih3ahuyOCSH2IN9wG40Ow6TIVDHbwlZzk9wtidRGOQpvh5YmEHlX
uKLOonhKv6jcK7iqvfqUKaaIzgrutVXVCch0MS0TuLBTniEoFw9A/+4JgymuivjjIklyL7Qu+CqR
qEec3X8YDLV0tDd3njubBGfeYNdKEn0qVmEjfGyi7TQdkGuY1+jBAyorRPJ8Jb8dmxAcZgjXkR+M
poO0eKhDl5NZaNly6z4Fw/aIWCPVnOL4g6fYREj5S7+7LtfA30ThLSatR5avam/vYwgVaDpDw4Es
P7E6QLFuh6XsAuz71tKl4t2/DGYfuaQ9luCw7qGs5EF/z5w0/5IPbeIlZnJRir1M7XS9PiQ3hkn0
3M2mci5JwFIvmwO4OTyTsc8K65fd6lNMi3ph+mPgW54nbOWKdeN7ruNFbrMgHXioCVJ1HyjvZyVE
nwDl2+WayhD01dciF3VtLHsfGoYQf9OJe8mxRH/KdE7beDcCD4lS2z7DIn0iS6CRgOIRafGLPwPG
o5RvJboVpCRxzYY4ih4HhufrFezo5VFcU0an5Hf0WxJt4XYG8sgtJ3ccEhxt7oxPqag/XqeAhoPa
KsxeISWnAqvg2cVmFzW5+TklX+/QHXcz7Y2tJfYAgbzNHQJpEnMkVtCf9NrMNrHSrd5l+mKbYzKm
L2celAk6lA9DT97gRFTYc5/MugjsYXQwau4fdtmuuLN+Zqm41ukqmU+QZJOI1yLTTZYnfDMJrvV9
+gQTajphzpCC7TOSRLgiepzacCr2jLljUHKfWKi1ufOvFCHDrDQ1CiU9u3y79Nb1kCzajmlErodx
bq5Bb2hIGX8cMlpsv5T2Dtv50d7FIGePTlwn+T8tzajeALHgI//dhnsxTbCPoFfaM0hoOIq8RoGE
d5NBpXPKh/in66hvh7/7YNFQ1o51Z1pMJoeJxIuayn5tOqU5JHDsFI5y6WxBzqnWpfejPkbIH2H5
jvFY6pxH3IyhMD2bm0bZuo5GahY5JAV9hRWb2vXJivYa8zZ2DubpkdMQ0jounEn3MbOeU5MPkVw8
fGZv7y3T3SId6HJ7DP0RD6jTNOMz6oS6aDa9KOuFNEnKGTfuH4OJClxJOndHOL2R8qwaYFq7WlIp
EVCJIV3yYSGGmnC9Rj0XuzUaD8yQNb0GmN+uYf7sBx3coIJ3EJpbu7i615W9o/EdWARrTNq2w1nT
8D1HcAMK1AVUTGQo/rVM+qSICWxjVFshjHoewGdJ3z4RFHva5SdFoliiMoqN2Uc60jarLQDWuhgl
Mm03d0nN65nZR5bbrx0CJ6/ysIGfBbVvkQhW1AwqIis1YjO+rA79fTrfKW+MvRDpo43VDZxrw45/
1f5i4pK0a5LAKa+ulePB/jQqWKtphWMBTbbY3tL42jYA+3CW91aDm0YWJmHxRRINVRAWCY4D7LdX
b4BNOAbk7fGFfjip2rLnja/vswhrIOdlYPVnwdgCdh4a24vIZiMwjrOvJJLJxRQQJnCYhXZxM7Km
gyI6X5C+DMnviXLP0tt57safkMhqmUgXGfGEdnGXXOYzXEbY4/FaoVwZuI5Inqlth2qTXtk6QZQ0
qJvXojCrHmusz/H5KLflLJ17JY7BHBW9bYNq92nlrVBOu3Wp4S7J92yosOPfHQ0+F9MRx14InxXd
GtDgMF+OYyXCZvP1jEyfwgAQkfQzMisYBgCXB+veybzL+fzH2svwexaoIUyP7bx6Z5ygb4Xj5jBf
VOM8pOHOgRhbRIFTA6pOWuuC+QWOBLVFEMtYYG+DxNd41KjJTcfJ+uA2I//htnpgoCoodOuJcikd
bL0yRz2Or9+0GrvKW+ojXNTCNNrW3a5k1YMHMqRTg7jwZ+dK44ZpOiXJNa17hy9fimghseLAh2qI
8CpJ9vbz2kqwxct+8dkARfH/bTTPE/81kb7LwWLxKqN9xIWs687SGfq4UFcExIpwNL//cR7Op5+A
/Q8Br5NRZkmqIScamk1qw341XVhB7tlUqgh1mYdysBy/c3TmOBUJYUuFrlkkX8qPAFxKve0wCeZh
XLHFXlA2A/aex9LkxbZWdWWvBBmv36hF0EJ7/rLReKj1JrMEYa/7SX16Cf+UHGXWmABTSoo1fhQC
gQdeDSq+RZQcEbwJ5CI+eQiQQQB1oq+RfV0hX5g8rRR341NCisDPlkwJ9Nxn6v/j/qiP+i1SBpgv
berV4SKXpu/4DlLHQwOZJY3bWfvS/1tTUh3c/rDOR2271a/2hJauG6YLfCYz2zpCwHS0dnGzPVlb
52Dgm0K2uCQwzZmJbJr6/popOY0sYja7ST42/AV84mswRF7OY59nl1g8QjzWt/3UguSFoeoZgp3s
1tREe7GEsoa8anYemzi17uHlj98l7LPW3nPe7g4z6Hx1dEEjJd6g+9qY9ujpPbENITvhZoGUTf+V
HOaeGg7U4uvU8FVogIR2DsVVa2e0QQyownia76j40aJEqmGb0/TDGwvNgQsY9frZ2YNhQjyYQfrv
z5gm21A7uXdXWuJX7DvBVmPMoNPRwon5txodRdpzaAAA302U/hTajc2aj+sbwbj1MWitk4dSE4xW
PJiOqj/O08x0Cs+CdYKuAdfGDFw/W1qiLGw0d2eIIoHsMtDJ52MJm4kv47ia+sM3HqHeyGIrypzr
gc3VZMGiWbLiAstkDBqI6Wr/Rv391IXUAHTJ8RXPxAYBEzVFkwZKvBQDC5NUfKYEBvb0s+6P05vM
8o4LKR1cyzAIV5EVOd+qGLjRsXR9l+l2R/SyZtjEpbdxaVKH0j3TvbupqbOaGuzvcqqw3cQcBb9v
cEDzLJZ95XlVMWLUUSN5bGMTDW5/+LaR9A88vxaO/5Dj6aHg09kFthQLzmmkQd99L1tmSC8DfseU
7CjSoV8UQ5sE2vtt7+yJMJTlLZRx7LOQ+asw10QouI9642PRm3yjMrJAbEfjxLhGmqWTp3A/PfSN
1WpwrXXdtvlsWgNTljMnKr7p8Sx3ExxnGQgeFzj06UC91XVoNodL4DdImWh1RMoEVn6zjA3kbwMa
QP4cSKZX3UA1pIBI22KXIDj7TWDAq2QXZv88gvHxeseajZd4L1dXRDiu7hj15sJruMkYN/LOWRe9
bG0M6HEDavuCFy/K2uj2R6gVYhs1bwuXXPAJEHlIZD0ZRDqmA/VFQQgldlkVIMrD1uWbKqBVYz72
Ptl89DXWQ1n1QVZ1vd0U9iDxkBAL2+V2A1lSmdZr2dVAcCWJobgyg0fI12nLH6cWaXvvIpBntCth
PRPTaRE6Ze+E0MeDRQsNVN4YbBTwpqpE3h3SfN+MwB7kO8FS41C8ie/6hWPHGv5AToD8GJxaszKH
tLI+6lqxBHYN3cGgEJW6821OtIEOw31m5dkawsblFdSYlEpA3U/QeVUhg/anapCaL2ahSRtyHLuL
UuRNl8IOahkPIvGfB7Xg7bLn+Njq9zlROz/x21Ly5XhbvEGmDx0hD7LOx+wAHav80gJcj0a8UUJT
ThKFGZD0YIm9GSw6Us7U4uuabCBna6ld1pxENEuOtAsifj2NWsLccPR6RkYcliEF5/U1P79zBUoO
b8jwn3SiObepab/iHqP2rQTWJDG1cQrfirKLeFtupPmey/X4h+cGtlWSn44F33qAzgKCav97P2Ve
t/fvA1vCMWngfHDtmXOAi04LhF8sp6/qQj+3Ecu9M6mDHEHmNHemXS3hcddt94VcFO/YHLOSnMLg
Jsb4y1XpiRuBh2FE4NL/d8+iQb1CGtWGX2MejtkswN+/IPasN4qfeiIL9VEoLFUIpBU1FBqXyOpN
jQXd3rfa6WvAAipv2yk0mmdA4gM6vI8sGdPJpBaj3R/+H4wHzz8f+/4WFBrZwkrw/PhYCuW2NAC7
Kyv5Dnsz0xT2+tB+04vDxONnPTvt8nwqpAe+VHXfiz9otHFrEBFwBIXPkz64crjjVTnqRWflqVLk
igpq1Qls1e0a1XLWBetGcMpU4ME7Id/19l9bn+BrpGWuxN4nm1fya/kG7oNVY0G7qqpU7+mXDTXw
e+GpQa8qS8Wpgafp9a7SS+WqIJknmjsVDM8IES5y6JZdL++tjQ0HkxtC/SPhiM+120x/hi3emCoR
jHgUAXTQl/8YFZS1YSR/Xppeh3ybsp4r/Y7J+rHoit+EUa26/cxErDGG3WwEJiglrTu6Vc6GMBbd
jnlyageBOBj2/ojkR95nop8eRHg+u7qHuKG40VqJZtUD87aoRLJZSqoi/amIxqoVgWyJtppIHVEn
31eEd1GcCI8juCeTkUtkRg1iDXtJVZgoZM+GZfEU2jPmZOR2qzJ5qTeLgPOdypBr/bZP6qGB84AL
WaluEHtEiKZhidbBZTmkZEUgXyQ5vZrLKMxj590+NbiFRN0vWaSLdOLAENb+ow3JG91CCZ11Cf9X
nsjH5Op0MsxI+fpBc0EzbE9j+Nrqiu6pzGCr2zRqrrejMWjzYNiD1xuNnE9tnzR+iMCbPh0nh59G
c0Q668hMqI3wIAf2sR6DxWMaajDBxQjWrrmwYuLm+a5pznMdh16o09C4MTKULGJ0zknhMLG6R+zt
sBQz+YJeTT6Xh0VITXuw83z06EEKnsgVUGTaRnGGvU4P5MR/+5dTFIvQaAHNjdhc+u2f/iqKtNRp
adIAngvk4KWAkGacbXGTMwkJ0/Ll37Ge3+VoYW6xhE9hJTihHXHK1jP9hkn+wajsz+2KFE5FNAs9
1nP/YDmbQnVueZ2ySJ7txYeHNp+iMnlDte3nypdElHbYj7FtHt2yQO+4orhjxNKt8a44XXW+Svey
FlI3+86+Q6HImxSj43/aje9SbE/Wt3AznNZsGhCuq+Eps0Gl1H1ac8E9v+XlzZ3LSyoybYm0UmAT
bxHF/h/Mycac0bjuHCDXBF4Mox8LjO6X4J+Mtb6u3zd0K2U5Qw4/PaqO9CCLearVg0W7AiqOj0yM
ucbQkWFoEve7SabF6pZf5G5LvumrrwUvJeouVqAxjNvqji5czuepa6O+xwoNcIAHzCDyJSzfM9xN
i9D1WX3/4AspVvayEmibpHYtaOPYS3QnX8XO/DroYTQL/20fSZT9vNK/nAbsU7DTCctwrjZiYmly
ypHg4UdixOnw2yQqDiLJ/moxpvkEeYzZcWnMU6iuX9hg0u0++hZ7sdtU5P6TsHI1evqR1D7cBl+8
oh9ILPk/SQlV8VJuEvRwBvarFFSoweTi6GYX1Q5Xh/tpR3IVxSWagSFrqK/f6ylloG7Ggx35AWb+
yvbRjs/6B2sbLHFbm7/S5MfH1PLWdM8QMPxXaLlRzsKiV6PsV8fnAEhCnatMCQcpFoHcAl0E1ZcC
PZx+i+vA7yW5CQEm9pygnR6m2QyLAfZdjbc30ZWXfk1eAQkCWvwnvmpB0b4bNsL1lzALepKRTCbA
eh9gmcM1MC04E0vsPKFm6qlRahcWHywILBTBhxwHS4TaJwAJsoqPueb3208Xe0TKz1JYfRmmJA5R
21A3qOz471nXhLBrE1hGkcMIW3tXTK3xkJKFDUxFWvNHuSfylfp2RtAAe3UXPn2fEQqyqrYYWRRG
3cOb/WnThgNURnjf2SU32Ube7Ur4B9v2hdYxnkSsiVVoGxewhj71C47iOjf3TK7e1LCS1q3cueFR
374e+CQWk2+rlWmwZZTpuDsU+8x1fTSSu4KSAi7k615264IOARj0oh6bjfCGpEJs3kSTWxAe8Y6O
LaTmQtzTi6iO3a/wXKQ7JNK2BXoPu74LzDoowZS/v3j3mxaNnZ7iuwEU4d37g6IUqJRwX1I/1Jpl
utLOiQQvN4kHyo/yYmEyL55Ar6kwBK5kg7bUtb0n68u139EVVeN3s6aolDRmuMsNBda6TUVFWy2e
FMIiqfgNv30iXwWGc5CqhRGfhVvTnA6A7YEtnwJOz+nvnz43T6fYW5OxpPHFMTbK0WOGN6GxbBKw
zJH63ziWVaDCCtmmyAjGyU0cJkUSo9iMBNPSh7v8EclT4Qp9YySQEV0hpgbW7v//g1iEa5Szg3aW
Cwc15kSiUwf3RBuJKBiW/0OPGuPFG0Zobu7zQhyrBF1CezMrxa4viYQQOWWLlinjx37/MNO8RfmD
NtVm7VND2qwlVcMDVi2qToUkWVV2vtdNugMPF0hamUV11iGjtBmE0CRmFu26EDiPV2Ca1MfF+Shj
IEt/uXuAuW0RKvpN7kkpxVEJv9bzsZl00g2O6PIoV55BTiA9lb/F0g1xjVnKjfIGtYzDNNn1tCe5
udzbeR/bmQ5LdtS/E8Zd+8qJU79XPA6z/n+6DEc2oj3PFXWMYgkCtaPPoxXNHSR4/77G9RnqcrqO
w9VVi3LmEZRYQq0VD38XziusUGnQMddzSJQp3BA0AkZryhV9kgUJsEQPmUSxAdQ5OD7c0nNpl6bh
JUYSfEMyBElQNFl9rza+QvCh35O48TkAxHLJY5ssdogRGFu1TUe3u5WRw/7Y4R9nAScjhXT1Sw/X
uwBryGI5NM9Nx5tv6bvVKz2GIGJRjfU6lnFVIv3KMDDCzNK9AbdM0Z/RUZygUV7gj8SqoPfMy0a6
zJXdUIy+vuJBztntUuYyx+mNNMf69cRoCUPEsgndxxTEixQgPoJfS8TGzb+NyMMvrD/yN4rxfPP0
WKZBxSo5X08/b2tLpzoen8dXnoktKbUu1dU2Ja7DD9HiAaiVNLTgDAak7cQW5+Ho1/PWk/ab74FD
/oSDLmm0vtHhPDjwYud4KEvKY/mzqlZSTGr8KVgnLNp17Be02OVj/AWPjWuTtEN0TTFB95ZUUpof
OcUGdw7JDyWcXkXIeyi55QFT9665Ntsgu/myDsTAV6hNPM8hJzErN86UlTX0uoV0TuVniUaIOxce
uNvnwQehqdr/SE66NA6sKWWcTj0a/v5zYUj+v1whrV4qZ9LfMi1JcDGmqbSB/ck5pdc/sqVC110q
Etb5bytYAFPUXdjYI5ImZ8FgLec7H6v80eoBQfYvRO5/9R8bJA/FdYLpMejpiY58W/a9Nlo7Dy5B
UiS1D89fv8Vvql8cS4GzRbRc2+JUJQB2G2xANMweEVcd3iSpXAnjpnOTqUFPiiGldSkNYKDBx8F+
iMzHkAZ6h1Gbm8bnxZLW+vcGuUbHaBgpEpV3n8MQskBq4cbBpcYZ+W/2atHq7Z2hhTD9lLvStSng
Q7GYDjA+Ifmoyr01EFe+3b9N6aipq2lpQFyQNA7OrOGLBgiUWEgZcKZgsKrpfSHih+Z5fOQbLVYi
wDmQkI8REQSlI6qO1Su7NqPzxKSUApt/R8Pl2qccJ8bQ3LYPFIT0kGp3En/ak1G0dFkvD+n/DdVX
J4oAno2613jrzUapIOPHm5BA1u8bFUzBVfNgDdcClRiKg5J+udrHlCYJZAaJYDWkcmeQbDzkjF1j
QItJuXF754NwuKO4mW/Xzw7MOUtOUk1YLHxQ8oDfz8pkNxhqs7VP6DwXh0DjUU15dlsNAn87Dhc9
fqXdfeHzG5c2zxFot7XsH7/hZZhVsdhLIK3T1Q0PzYtlez1yf8rIZHGHrbgY2JZkJkIBe/M3ZGzN
PPL9V+L999cNHbqNzStxZZFtZewoa/tySlFlgwLfQDTpEZazADljA5saTK16IcWyMlmyRRaKa35o
pdv/0hLZh6FuwxFKKAqBChE2375K2ZCmEy1Q4Z/oBKr8AGLTjZcBXe7UwfST5W/4oNaiYX5etoPv
OP3VoVuLvx8ZpsKrl8bAQ5Br8KaPSCsd6A59KFvNVVW/LibVw4FAHcC1J3z7hf2myd4lxqxtCLJu
4kiskoO5ZpRrVyj7IAbdy9BF7EWFDJCNsGm2ZOu8RWYnL6s+WFMzXZ/TPGFxgdy4hW9G9IziYZh3
9QgO+elA0P9/Xin7t/VkiDSCJfvNP1tNI33VCrXizqAlrn7628p0qa7zoRsR6kvqOOAiPyG2y+9f
CcKP4MhUVJXdCTyh247VDlf9nBUdxf7aFJJnNveqTVMJL0P8Uuk35G+yH4WIGw7K2jx/biNlc27q
EGKtbpRV/KotUOOm/4CUtuo6WdW54pz1dAfTXUMYGNK8fvc10zUJqWjqyeRG/iOPIB2hae2sw8RG
KluY9HijiKI2Pf1E2F60VkZ6JrxhVETEcXBef2NXEskoFEMoyppHo/YuEkO2PqQygYCt94XIyd3c
580mBPNxw/wmSxWMFIhmzrm067BjeOP5GSu+EfEGUGAkdk207rYoWzFAg+QvKqKrTbcPNgnmRnn5
ItnOu54UzJSzQDbMtjyrSC4f69hdIqXOhU2dbYlUJE9WXP1p+ROQagxRAs7UT7jybyIf5zdEQ14E
X3wDoGpTlTI8DBNUspwxOVB6eGCUIBY2X/VncRANsLf1uaaUhj5/zlccBjkgm4ZyfXTv6wNSkpwB
OWogLG62sdZsjQ1T80UjtSOOGqgNZSqbcJACOlN1jLN8VLi26lRoAJDgcQQJPUgUlWsQNfSWfODu
mWdiWKRBL9+H1IN03xIFWspnR5Y1jsHGvskjNYS3lU8j5in6xFcKwgc3cxATGJ+o/xARDEM7YUlv
aKyB1+CWyUwOnjbZ4Wng3ncTCXEXjZszSiYwOpNwDsSxqk3wSLt02ogq8MlB6McoTH2pKmC7+r4I
locviDwh+QEiMJRLGN3xt8qtFBxV6anHp+u6HHptfOuigsNydW5lxawLIdKelV24wbqWGBQEk3zP
PdRF+4vx0PygIc1jsRYt7MDQD7bqxVxgrvrbqND+7mwxtvAba0bAdH7DMb9ksdcYEbv7aTc/KycB
rfcgLHbfxqalQBLly+yWqrvNIAK6yOW68QIK1TIEmR/9mqOU1bCojr1BRNyfUAMMHCKJU1h+nAE+
VU9I0ocY6y8BqBMWYZC0Bn7aAVyUO7w+N/iEbGC5d94uHXRqJP9me7vDp7t/gor+QgMCfRCrHahl
vUJfPlrw9aUo+qBdx9NExW+rJ1o2S7x3QaxHh91wWBO5biZDN9iXWNW6Edw62l8jc0vNh5Fqbl5e
1mg4UICzlm0aPvwXApOG6dDMTnMho8kOYoKJmBnYLI/oDJQa1Y/5doe7yoWgO5nUSnmqw4zfHZwY
1+4D3MBHJrvo6/mcdGLqZT0WLOHRoFGdNRDz57eF6aIlyVMGJhghggRJhyVP+laav18Xckqh0qE2
Ep237+0fmCbC1I7cq6E8kuk4a4A48MA/VQVsgvcuaL0tOM5lOk+/qzN4hMtGqVktzPlTV3Mkw3DU
jtQ96FKYzVu0nPahliJFdF4FJIufjTjbxEq20/U8+RPeg+9WoaT5f+wycTMagDZDN805dLlwftIW
su6/W82rxMb5rhrEwCOJgfQF+6lUWMWZen0caeX2pkWbjZ47ovPRFK11v/rOZzD7xiirvE/iko2L
2ppxTrBO5F9/XK7IgqfxYRb6bqV0k2rBoHiXTcD3uyoF0seHJqgbp5uDHIOhkxjdD3QW2wF0u2oW
37TERVn2pGvAuMB1yUCWcuTzd/Yd5iafY62THe/ReWIyTUXDuTYwUh3A1UTxQ/O5fUyJbc9delCm
SIeihL9J3RpoiMy2Pi2hjcvnkAY+3abGB8vrcVvxloGaZJ0X9xv4DSIoetwWwpNCGz/AmQ+r/cte
glMte73OtFJmYvbNfnsNf/nmyKA2+Q5w1ZNCAvty29piBJEdcsq7OpNS2dmcwv1qxBm7GaeMU4bn
FwTBKpuYtgpxUsm0RcgNx7nZ2WGF0wHcV8UqhVUE+BnfBlnQ6ItT+2R9/b1eMLQn9twU7iuTSZLy
pyOyXlleEyxDJogKrT8Xv2CpTletLIn8uDaQ7IQqOi4TdpCnMCz5kFom91JeH0Xc3u9D1Sn9+VPR
40XgEKErs6Y8s+0PpsoF+NIBWOFBvN48pcLOW4UgIv0teRCVmSxi/zteYqm45Y/mECq7Fcxx4gUt
hxtY8ar8K4/YGAnnCLhnYhVsIAnt5y65nDEO001duAvQs1al2Rl52q4w7vkORKC8VJfb/ReaGo0E
+pfBEwg8x0D0sXFry2xtcb/GxJN9rCIUzY54V9WhllwDS/INcCHF3kdk05EjtsAqLk+ngr/i+wlA
fAiLeX2sYAGqyW2Jjk77DT9sK0fIEacg9d1y8RqKohZebEk3o8oGBu9Y6H4kNpV7jFNjvjanOyvH
m+QuwoTqTB+x7Ki3eI3bW3JC4hxUB3RPSulE4znM5/nX+G4XKg8a5nQ75jK0xYHIod20cmCZvi6c
hyQWvvNDWnSKiFclI33qAL6JM+GMFQt5CMtsYS6v5IVyakGp3e6DHsYBV4knCy3CRAvbUN8dNPgE
R+1iERMCP+27RZWIltAd90qoeKUDOzFeqYHiWw0ie0rP2OofTn9RSuNRrEKU3v8GlUafQaInOeHc
37OgHZJST6S2HPI0VsyS4yUacOtULkjpKa/blujdoGuY8n3mizCwDGXGrmYAyLkDhwy97BKp0f1P
TV6gecSLW2iReH2drWiLNq5TIZuIJ8pJ/MPe6XInToZPhRUuXqPAUq8HLG7ojwTW7diY7OD587UJ
wkr1CJu5M8N9jnsgsVikZdzF0I2Q9mrDPA9Fc4CsazsifeakJbtmR9RhS5R1bwo0LFeJlp6h0E4W
psU0O5FHk3TQMcgDWXX4GP/2qLUY3Mm7+dcs47zb67AIYI3dFu4OPgVRQgEVM74117Fr5uNp15Xg
Sj+eliKMIYeAW/IeIiHDtRPSRR48Bkiht8ki2ltoTz3GCWmtAoRx+bpwibGikjipjBWCI3X6c1Eu
Oh5SYfRN0Piy8PYb9MDTyPe81wcFzNd06wExtFhISE7d1tFQDxGKd/ZCVskvT+Xpegk7eMufHmZD
XXJf4qmMLQXAfRZFEiiPndl5ZsfXsrbVTxUa67bnCWGhKsB/UCRTgOZ1PsGTKvaUAY3P2o/lXre9
t5pYVCmQkyQ6HKH71sm1whyjsD0xklkrniyzboN2kWH4HnGEa40vPg31N+IcFFwNzU9Fi6drtovW
8WZL4YyyGWestPNbEY0bmGAT14OhAt3kyMi7UoHhKQfT1bc285slvmNCTK1A7wN3ISYvfxBms5M+
zcN1rQSWY1j+Rkffm7zALfACgM2DdidZGfbvIvSYvqxMtCJfgEkEdoC57T6c9K7iFpPuatOfXFL6
jGDEipSdnhXErw6QR2FOOKM//aObiwTgRdD/gPucfHP3viVyBSceu2cohVoxtlbmAfOOC7pPa9Ii
2sf0YMhncEnXYZevD5oK4dnTt8Gvu+FRs/5dggJVOq7JhvIu8rpXaIgqOcyo3tPDENX30gk2/3aP
vcV091hRGYsmZLBn8RAeAE6dNPNALFq65TMS0MflHiL5GFVceyrD+lr2u3aQmmzuZ0TlN3mUScOZ
/tT0Ka/5B0HBSPbSyV4g/M7HjG4Q96KZmh8SR0oPtGcjnJjMB0r0stMa8rd0IEwRQgrfjYi0R5aJ
s4MHuKpuoqDm+SJxQNz6ELkp3hnu83bB0P3BeHWGnUtsJhcqpmoK2j6+dXFWXHD/+DywfaWbchE3
2Rfd6K9IwFIW9H2TwXml0LeqptQ8xErt1LeR5yrmflflXXT0muZCsrG+qKcOc7IQlM2qYmLNrmzP
84IK+Kbw9TFjY/dGhE79bu/lFRffcgFLPdMwPmt+IvzEDX7L11NE3ADQxcpPQ00Gj13zjkHV8DSW
uesBSTSwfqDZ+V2TZVumv+MuAbxHNOXcBxqrgy2fKEDzvDEiDfZjNqFEXPLgN6aOeRoj3ppnl6nA
5/KaJI0jpsjP9mICMzI8xjmqIWx74BhwqKLRbHWSIGFzYJ+V+OoufiNgwM5X/HDmV5EtiiBUmjL+
2xjvp7Nu9ObIiEoJyI5Ed8KL4LxXO9u+hOUEXpgboiU3Xqhlb9hCSGCclWkajDSic+dI3VjrmKny
YuzUsVzVB8WOqIjL8L9RGZ/S/YM4vKlhtLCs5Oak2cu1SMUGYl9DyMj+ZXeKE7g1+5yZKvCpAuyt
u6kywD9K3rgHUKQXS+DjK2nppeZgLKZ09sDpgBY3ZnkYrG/7lvn7n4tSEGWEpAFNM7AMSNkC65dC
BrX0LCdzOkcjuAoLx+AXGkpRGr3rfK7WT1dIa0taLe/BihTFEqO7bouD92odjmUsG23f+rEpK2gh
8rb/39slwOsezeGfKf1FbjIzKKCX8tcyFbH++CY8dqlbtAqgLskrP+YX7KZYHfzhxX0AawD4v86C
xJkdJs7h0/DoNhJ4jq/S0ozbgnkazavVyy3hrFcAxnSaNEOowRUgmNAh9RAYycdTdbMnQfrVMXwK
sgLvNbfMJWrOSLOESkyOt68vHhhO94ff4Oi46CENyTTIKkFLufm8gj/APlhaSGZej08pfi22AAXn
6JTSOwhg0D8a3ASOSuLacyKoUbANLBVmnyJ2LkFGizMGBU6e73xB3SaIafEMcN5bRdmJ32e/3Xlk
JNRwtt6NVc0n3z0IFrWzVTl6skD7RW8f2Q8G3Rvwy83RWyja1k6a7QJEHi6VZcYHDrEFU6Tltcmr
JnB1QvSve+FljZxs1dg/xi5nU6btrHRJhPVmf3Kz61DqpH/hzadJaAngwmhU4B8vKfSjAzipSByV
0Bw1ZpdITTWdiE4MZE6qgk7nMcIS575QdSb/bUVFxfPqZc2U2vImsGh1bfEeC/8brmMLS0fzQYqb
UEJhWHG/TPOeG0Hcu78NMJnA1MQKX1UE+pr6R0KbxsI4/2syvHqE9YeFohIAStMZLTB/T78HRXRF
AS6/Ix/9ZR6i3Bjdvg6ATj387K1btmx2q5ba2sDZtIgBGzU+m/RB1acWr3HkSSP7ozoSnGbzBq+W
oeD/S7xFxp/9ewVl12DMjCYMw79ZuG+AJA5SfLpoOeeTH2v1Bjgpp85oKxvTto6CA2Bl0PhWEvSK
tU/4PKequy4vOxMK+gZg4rik0kjWqIEQ3Eyh1xYhEy2DTDd3cBa2A2WfN1TzmLPzNQunvrkVh4lD
0COomNr0EmIHSXaj/Iu+eOQwQ3EFqLwOy7fJiKfRFaHYohYsaZXCYefpfhGCjui+P1SgUg5tsloH
2rD1KbC4qG58PzFBUzBIw44iQd2JxjeC+cRxaWi3YLL4V0YYPU1qkGJ9aYFA/LzQQZ/ZopEdnJPz
iJfn/6lLmdUcfUtsxD6jOq1ZLnzCWNT7AKgYrDLBz9vTknzMIPprdQgTwYOdRnEv4R2nUZYJI/Ha
7OxdUFsIOSVbU5c3IGG8KeotYV7MV91OkkdIkG8k9HpHFu7WhUWqrse2D3VXMUMDJDDYCTzLcTOX
FwN5lo65crX7NU3U/kjSiSEa9VOZYjnTsB34rMSA4MXFrhs/go+be/jXALdhyimAxS/GHNjIlDVd
JmkWkQZx9F0LV3WWNhk+Dr71JhKBph1btP0aKyENx9RBtmf4dU9MU/J6HFUXc0jMIp0PP5QhMgVQ
4PEdCDM9pvGaRIYqqdOu/Q52UlHW5lijBzfcJDgLqseyBGo84K34ftms/i8bqOwBNQsU4B+xGxge
RRod35ZFN8go2T94HNwZkS+MqXYCWVc2HgC4QQTew9GKDX6hucRah0os9hZd89XBHrtD9GfJqNdN
vginVCuUgu5qFJWzOvCcAF9hveBLoa27IBJO3pausFbsa+k8X0YPkh6kA2l+357i6rvl/lg1TFK3
sUZKFvrYFSA8SFkkiS66vQFw5X5xrUJh+c6xHeMtfs7GVsahiN9kjC6LimqNSIwVXqPzWrcewMt2
A7Pfhgfc05sxZfMRsnPfSqin+CXgcorHNAOe3wyPA0vJCvEtoLMANHwEoLkGYObTzPTrGKx29I0n
cw7Xx+E7Q0V8IrciXLXmy+vVS+O1j81ztv4j/afmevoiAYSm1INdljpMMVmOpvwOG9/dK2ElYUtA
dJwO8Nrg00V7g3H+DmQANuHSC+k3bsE9QLUMwgxeCVyh92c9vqdz45/wQgwSq/C4fZ8P+fzp2hdR
iL7DtpEo0fgMV5GGhpwodOpX3EMDtklq8vHgRnlblgwMYEcNIxHs46YyKwClhACVEeJe3Wflnmtp
D0QGCAn5iyvdGXZmw3Q30ibFqs2+2cfEET89e8UJyTlwqtaYfE/prTW0kwr7LaPCQW1Yb0HfMrf8
QFhkdRkG5gMwUAhErDZ1Ro1zxui3vb+//pVM+Aox8BhZPOlckugLcq7D3igSc0UqjvxjSXaLKS3B
8K8PFTQhY7LdITrY9JUBTGRWx4lmBpLAubrp2kmtH6+Vy7rFv43I4POKKDLIUB+CenzLlHbKc1yK
iDz6nCHXrWLKdnC4LqdxfL4xt/4UzXpZ3TR4HIGCN47sJCq/0sNOyRN4z8NBD57LlqQPRVOojSy8
XJu5FKboC8Z2/NgTj4bGaMTIVXPUsHxljIfueLcCvMulpW8PqoBRX67aD0kRNkNKNBxFhl+H8cRG
FhqBVsSza+3cH6vsPKA7XPYR/O+GmT+k+sQHoKKqgZYdipLCywlNpedzZwHK/2doixG4ghtf8hVO
Xcw0M7oAuEWa3ef8Gqq8aRNxhM/wKkrEvHiYcLzVoJVHcJxmw3/s7okAN4YqP1kN7m2wFeMjk+u8
gwfN9CAK1lXh/Txl3+nZneSnqj+6z+d7kbmAwk/8I/11ArjRTlEFNkF/URt9fkEjZuWOSHK2ybyh
+nGCuj3BBHritbFhCicRS2aM+YQyifzfpp9zvA9hMd5Azx2GnQrULnrjkgapxvUBVlkVZBMuVRmB
Hc2ibeUqZA4xicIoZbBHhHFB/GKRdSOoCiH1a9HqRlrhOETemeEF6HF7RPVQ2OChCZ1fa8isIHrq
a+uryIQPTkc1TusM+vdEqIo07V60bi2nRwTpSnqKIkZm6xIxZ2ixRol7xATT1iGCrSBdSqidXWWV
r/9QYWLA7tLpKvwt5qmNLMgwBuav30169MsTP7AhWiLGtqcj7xjdFYslvhxYP1NT7lFQJPb4QD3z
I+bviVAtx8SbolZ2OycJFgx6aapoJuQGB2fn31ohInL0dzekjtgW87EoC5ZIZaWCXbnMJTCpTu0w
RuvmK7t/oSz8tw9hQdYcTVEgH1QyyO9CwW4F0+O+xERvoFe6VHF9C0E5hdY85KbgnuOnPXo+n+5b
T3VKDge2qZ2Xp+o5GMahH0HnNnt9j4HRka+o4lWChKC2JFPekaVT7ak0ZuiXImrUddQICENVUtBs
8FD7EwYvnFwG36usHk6cqvS0j+3+n+PHc5NET1X8OeK+URJBLjxCxRb3go30DZPWo8SZiY8xHiRz
UnIAecBcI2XZrxO/ZsiLIF63lu3BC4hjqYsJuqGSnv51/WtjjSfZKsxMhdKcJfMWScsyRVTx2gVQ
FbXE1cRfZjxoH5R/I4o07wZ3ctb4n1vbBw7BYSPeHSXSo/wUnF00gy9OARn0RKDsvsnF9AHq55Dq
6PvTxVIMff+8YSORSMSGzyFRchLT4OAkYZMQzGZ0gSd9CRb/8MpvWHc68awbbDIko9uUTKzA74K6
FFH4lPi2THFxU+ARWzDGhpBnDVLuuRGScjty3T01zd9nYKAXZodDEMwaSVSGPWYQkAXf4cLdjoHC
SM5rjOARkdsnhxThvcBzvZv7aeH1NJmznreQZfNrDYvx2YGxo675l8N9zZ0CzYVM3LhMToSRap8P
bi0IzE4JdnYy0q+PauADrcZ5xCnBCRsDpsNbr7KMAg9SttOzY/KqyE1HAlV83TrA5maJ05K1guW5
pW/xvqO4cZUTY5r6qQTrx/l5Ziu/RqO3vSOL2vV9OZhjk85T7TCObLZXjPcnQW7MPpDomO+SryfY
MlPwm7wq9YG2EoToGODmw56HTbv+UvJCTyhBds0PeuS36useGHXRrZlnHiv0MNjKooLaFAzdbB4t
7e5lL5/ujHUvhU15mXdB869TF3tSddV1LSSMleaMfIEthW/GKLgplYz6e9dsNhFGWC1358FJNKzt
fzJvdXjU5u07cS3ru0b+OW4fUKy5jkS7c2i05uPMVScma0YC+hgoMcSScv9U2iaS+bQNfPnlXdf0
Tj8awnzLMXap1YwYlB+WE9raPq3iV/MUK5GKtZkIR9FGzABX3t9As/dlsTou3jqf1GVuyChsO1yN
rnH6kT1QqEnXtb8IwTePG9BfjbCSAxqzM2jEWQ39QYV/sGlrlxK1bBRarLQGOtTfcpFUwPFNi9iy
agQKw2RGSu7N8BxDw9rw8QdPx/8keCf7ShuRhpyiqPXnzDKyRb+8c1J20naPmahe039sOl0MuGW0
DKwj51BGS9VssPn2zexRLvYUPKR+ztBEbZ85hZq6bykA2OP6+8vEqPFDzkrdLAwaGUAlxbUNVYAa
LOMRyTqxWAEM+WnwuY4sY7JN3JfXHtfaUG8dAItlAxdr9tozCC3aAdKPb/Pq5aXHztS8amp0dycy
YX8d7NDDGmlT4k1GbNb2gWZEImM0wBhOpoOuEl/XYH+AoigO47G8VFJEC34Ncg1Qokptz1dlYdRx
PxM6/3fuOHa4k2jwGch3BOOmLIul85Dc3hENlGpfOpkpamrv6NMdXoMbuWgI3mrKXuIvw3sHtWnV
vdl+Ys+b/0obOBabAX1z+69nzSSUKdE8l5t0LPtaXOhDvIfmDJee6zRhnrRgUy/9VBz8SvWPruKF
B43jPN8jtEBtGdU225n2oVnuAjdjOHsMJAA+5pDk16E4xN/s5wuWemPAnL/HOPnZgxI6T1iPpjRw
89uyS3fDhCAMABb7UMzwh6Uw5l/LKG0AihBfPZ1Cn7YFrBD5ZLzC70kdn7e+rRRBjaOJPJXY8AqP
f44qO26aDyM5mZNI03/DbNWEIcRs7nwdGOXdGjQTp3m1W5hWhF7K5+OdOaawr4S92E2+akPcqulC
sBupm+nDAFsceKVUOYa6klBCB1mcM/Y2cwcnk1anzoPxDK1ZFb1j24gu1hZyIzqMWJVGzg/DPiij
GhckZITiyhl346j5NLYzo74RFZuxAV+pmBZA3J/nEewhk3pwzZw83lxC/yUN5QrP/pcwKDAKxz1W
QCly+9l/GRsZxD8nvlZek36i3C0MvkjFeye6/YAKULUNPSbO7Zg2MmEfOUc1Bx6eg+UeDHCvhWUq
1oLJdCefriW+u1tOW+URT0e92u04TNjjnzBQzzQBYAVIovTSSPxlFBKCHsXfKqnzHRLfUyjQbyBW
tnJ+jWwY7BcJWf3jFyfMQZ1HR/VSEZWLWrSn00aVVK1MCo3syO7ntLjAm48307z0RRvC3FyxhnLD
VUmm88vtLYm/Rx8WfSkt/Tyb/p7VgvA51C5OZa6jd7vDS1rAGKwWXRrwUHCbhEGkfzA6hqifITWf
avueioKrVWqfSR998VLVtcBu6Ox3nmcMhMINrond22ldH9kLkcgUtd70HX3jWltNCoVMhgvS+J5G
zk81HWAp39FVEI88M61zXd6NcuNnLZE38/TYkKt6Nr0jKxzs88HqfTxN/Go9SMlYQvEAj7C001fp
/uBmcg8CKE/LZorvgiotWhrWGOc2p+okLNQI/eqtmcaGcFK6405MtsgJoDHfWUKUHW/uej6WhEYh
6LfA8FBpT16MJKBg6XcYhbUUgH1YTvLuhw7VW8m/a2TwyaaX8XF4GtBpqysnzOE6Q0tN0apLgvwK
cw4BfiWelhkhY5DvUqRH+GiU84CEKbzQgx5Qcw7BUyTKX7/AlBhj31vAHodYhzzose+4sM6JhnYU
45YGYcLqA/ETOZcsonSxIArOVOmD47x9FxCiS1THKgUtei+ZyYJ0YYh+UIWkwRUuxP6/3Ysv92YC
opYUKZLx+HQAH5ZzKDnU/XRidRI5wWEcOpM/5HEmIVAXZSdGIzfj25Prg8EjSSjGAmgbRbCiV3cy
fXE03sF/BOD/J4iiHN3VNrUk8qy1Fz3pJZXlvA9NpW7zHRtKhQl4VeV4vs0nUNfcGxqmwJTC2SOZ
QXHsdv2xArDwEaqJAh67zH7XX6ff1Ae6FUFOd9Jf4DxRyNFg/bna026YgNYSJzNT0uyducTK/hLz
Jb5W7X19Jo96O/atJP10xr4MuISIw2i3vgUngc3bhun1ZIMizbqfB/py2MY8wJ6uc44y3Sl8VsJf
Uj4e2J8DXoUWM72PUvhDK3pF+ndl8lJ7or11r1elBipFnPmPBCYEuWrcYib+3CoQ0WqRU700nOQh
GL2XknPFy8WZp+1BCB4Dw0cdh3+kCYNBCVdQOMQ3XtNnNP9zqS+WvAaL4nWnZXsiQTWwttm14Bk/
Y2ktmBx73owWF32FoOYD6QNZUdPj/sa1h1RZ7Dga5FmXkmTV7LOMCrI1fJnsRFQDSwV4GBh00ziD
K9ZQB+zh5KgFGc7GBV5bM+ZvX80zRJAJlwUs/n83XFK4YLPMbBTJTH1i0WK2RhOM9TdZk20Fbnnh
5s5f9Sz9allwg4N4UMvMaXS7KrHJZUyVqu+XnKN7dHn7NzLHd8zcNpfPlnaG53JvJp0AoskG48W+
YhDF8WG21iVNenKGvbPXNKnxsS2FH8TDnZ7R8Fl6xEBzTR00b++7s4enZ0Uwfe0ILh3iAXM/znih
UAZtf2h8ljWbg/l6bXim89gQQv+GobLjo/o77olwgch+xC6z+XIX2o64ag2EFxyGhYbH4xPu9A2a
s0u4oLUWxdQvSMZt/oW2jO6rb3ICM5D2YbBAS2bh3Wr4oOOdFZjgUQZqKlD1+b7rpFq2SPMUN4CJ
/4cFel0tooPTVQeQR4iO9EfpzziDlVUh9MILJFcc8zZLMGXUwWhd2vhDSS/b9MKui8ExslDGSJFN
g/jKGOBfCw039hxyXow8KB25RKH3ebxaodlstddNb5BV51JVbLYW+JZ2nNiV0UrgmcERVb6uBdD2
LBe7cBs7SQzC3BSVH//g/aDhrcG8bkKNky0B2R6ECbupNa8M53h7NtxJ4ygLSSkJF8XHfGdntvUB
4+suCf23YLEviwl9k0+h3vY2xsTEqNEwGZBw/GgWak4ntsDdZrnMVr0mTy4IQ/vMIlWMrAyMHkvN
3gFtOFDE0lZaJDAAlbgDM2NWM5/IMPOhhdyPNBZWHAET2hZuIFrNgFB1RjDXNOpooNDgZroWzGHG
1c9wjSaRt4Fzlt/xi+8uZxEpen+rHZKGONbeGLYcOXdb29PRxscZd+dLmJgUNe9Qjz9KIn4ycYfF
NjDY0mI1ZGhZ3wNsB7eT/0V0HzmRmftAPgWw4khrz5MdE9Jk2DHZYANEAx8QAA60319aWYTKKW3e
qa3sVnbmpD4PeJ0C5Ha36x/qdqe7hH3BMhU6aFqrR4TY/TZHY3aUnn4v1fiZLBMJA5fnUqhXc7jM
NBX8mgVufk6iBWpPcbUVuLv4GWpmlJ0C1D8mPDImEaYlUyOgJq8WkU/kgEjH4kLJf1mwEznRXS9y
9ghqlaJzZ2bkODAOgF4WgQiqCTOLYJKuKoVvGQRHzCblXwvNQD8y4/NZTaFEYuo3tB3SBs7S6e25
K8k32lGUxrmteWpy2bEuY3yhs1PzFvGh3jy5xpJ7/gKGP+2cIeC5LBMbRX/BMUhPwgdCCtoTskd0
hHG5LmdcD9F43E27NnSkDtp1dten3gIUx8EWxJ1IrVn5+j+ZaQQanwQpoNeUpy0/VCy/MS7kruZ3
JXQ63XPkVGnfWyxM4cMIdM1La8WlITEiB4Q4H2eGHHUR+rMCHwFqg9k2Hd+O49esyzs4wCDDNpfM
W1a5YBgbtb0eljHNw7jlMp/0MVmqJLj6ZrLW9cYjPcYaYM9t95xhj9fepjID8Xs2lllug8cptJ7F
bkNk0ptX9DnXyIS8Y6hWngTAkGfOliY02o+OwfWFHrjrzcVkKkTklGHGYVpXFEY5TGHnI5mhCbto
CHCGRV78oUfutCxMky7femKtHDPVTPTLYm7wQXHXItv/T153gWuNUu0Ha5fO0k6rGz6A5QxNcX1g
Aid1PBhXTq0j4/xKalfrfuy0z9ZDdXyEvSugufRuGukOQ5b9rkTrXw/0rBRlNiBVbJyeTt8GKAWa
O36o2HzonRXn7+9oPiVW63Up/Up7ICcNLVRBnM75co0tS/OJRIeYMI+6HknZa39icpzv35MDIXYX
+/lFvPOQj8gT7mA/h2Jw5fHn6OQwqBzfCMTbJKr0H706eR6yEvjY4ozkfDCMCaRUcFFqaWtwVSRS
dda7tONWr9oPm7fg8B9VW51eVpFg12q1Daq9ZI6VL2xhuCcMAeJ9+ihFlX/T5b5b2sr/9tYJQYd8
tiTD/Me7u5cOTJ03gUh4YPUiNZdN+KyzKx2rYN/xOxwlU12KKbI53kQBbApKsiDc9nPQoauYiOe6
cZu9yTgAmoCsmd+m8Qo6qaQosbYlpUK1+U7UasQwgr41sUk5EdUEdWX0jc38Kozxbagov6+/92mU
h/T/1vPTPkS0IqpvotmnF9zUK1ovaA40VWocqEIM3AibRxrjYYr+9oOEAGdB0b3pHNfaPVyarBgq
ZnOCINcAr7fJLQg1dP1MFv4Llr0sIkNUqHV1RLVbJ8zaMsIEFIpk6mJTxkxMdAN2Xk241LXIXx+C
FNDWgJ5Iu1dmNHFijEZvI0CoadpnIItcJQOPLI0fdue3rNILMntHZFOELoHUQ5JmU5nWIxoV05p6
sLL1PRteD794Tbimu0JWIeN6omrY0tM/7zUgB4VYr32P5RvkUgEeSgXChC/uGP85T5n5zjZpTUjE
vHuYdNej6oXIQtqurwFLgK3heYx772ezO7Y3BFoqKJElOqwjU4Ibn8nlFVJb/9HivBlKJZA5NsPZ
eC1JU8LdB+Kx8AbuCkuCqu/Vo9Ij9o4Ve2auMLt7hCXA4+DqZu+5HU+3rgrhiMc0q8hLtzkBZbQb
qZjBaJE60jSGE47w0XgkdZknmr1dCgSR/7q3hXP1JYFc+dNyxibSIg5uSF9wVptldbhSeUoh8X1m
qBlK/aPxRCsVGaixV0r3nqXaizkHX4rODSI00VH5r6MW+IbtX2woe5uY8peNtBKnjJLKAhk2kNkg
UZu0QiSkfufRXC5Lc4FCv56Qfob4Ibusc38+cFhDIkse/hA97DSxToVqKlJdKxX9tVsGuguNuj0E
tdzrNYltygLunh1R+coMi6+pgM+7AhFUxRyG6O3rljtyJkIXveJ/wDNTfezX55UA1riWxVlsNTXz
73N97VLbDuFIfFzl2Lk4mxTy44ZbPv4A2+s/GeLBsK01tvY8pvgbrYASFnOBjNH+uMe+27RsEqMH
lPhqq+Q2avYf2UnPJg+XrrdXO/0wqZqoMJh1j5ydim+5bkLagROvz6JE4Q1PGtYqT/vXzUx5AZB+
diAYpGJsXN1HmUNq040b6YMjLupmm884K4UkA76UkBj7rIvigGE+7viIMtSedG1Q0lGdMOgvyB5P
GokKj4i36qJ8+vbt9lbaVwNydhaM6xHxMnT52YpsKmW6pRyZQ/bnYNQUTv+ctbr9Mi5kEPGUg8OQ
uFJwmikhhiCSMhgjSywegMbPvXMYgCsnUcraczVBrZeKYYt+KgbmTjcd4DXqmSVw+iBsXQ/muusD
WZAkBHKRvseXL3wi1ZsXvux6HqzlsV7R4KKjKr3r35+uBeEJCQXkKq1jMc/UvDczFZeRBQUFa/H2
UlNFaT4d327NW+tMvxUGqd/cpZA9Ag6F4TLTjXUcnMkmIgY9y9DhS5gQhbPbd4zddnu7GpD+0CH+
pTamScOwQ18bf+LkSwVS7nqcXqDaDQ/3ZAnerl1JPnnZrigWNGlm3QrGZR3xCzQXUGhE+1j/Fq61
N/y682e/jRrh5jBEuLIQy1TjJYaCqwzUlYq3PT1xUT3kRAP1oJJDJ1ayYO8p9vPMylceNoOIujGc
bP42ctC7+lNaKEHO0yAc5THapu2OK1zB/x6F3WjQ6wFzeHN+mN44+JuccSOjLt0MwQqJoLqNo0br
yer6rey04enbYTJ4Cy3o62fpJKlroEQOcPkyFu/13feGQvfNIC7GnrjWtbybVgoOf5CeNeE/ySjQ
+SVqm17h9LZHzw7EGYPh7xlt9vatOtn0F7FNB8ajg2oDaGCSR7lGAXBiL7u9hIrzcaG3ro/zxWI5
soA/pB+/fdyQD9Hn7bXGL9YMFzOtoO7kHLfuS/ZjT2wWQRVy96wI51GA8JSveFWZiBBE2IniCtbf
MY46JMY5j4RCEV8s1rFwcSHlbui1sX+oq4pT8bnUBSt2cGDvjve8m+SvjDuoVfYeoDFFSc9q/Kl2
rjUpspYCPj7L7L82pUEW6VDeiOa8SPvkGo/ksX4xLV9XhIhPubxrKqJvowIuehSqp6hggWhlFEcD
ZMLO9y13DaROel95jBHR9Wk9wSPSHBN5d4ooWQXYYQnkb7MSFi2liMrLwI5kpTXgOiOZOhrq+WK7
RhWiq/g4VFlChoiKHEeYRqSL9hDm3SEkp6Z17Nz+BgHTV/gM7xPFhCvirQ8jmM4HJWH6zn62jLQw
1nUvPHo6W9VAcLQIfl1GTClx5k1nmJlwLnwHCyEUixWOR2idReAnGo8jhm/t1hMVN3P0AUScen9E
dr1QbsWiqt3vBxAhX/DuGY0cIIhkynThKGXGIU4urbMz9+8gPsKF9YB5QV6feMYiV5yr314TcRSa
WbaNh6o7pp80TnSXxfgEDk/ZGW9sXAv5PYZXYks1usWmy6gOHRDSq9UWFEycSZIbM86nE/oslqDA
4AboEEMi/agYWM2btAoGp2TyfwKLH0ISVZ6itgNP8e+MVv4HEM/cAK0orWGvKnBJ2Lg9YB4YUZOz
32rz1j2oJumroqHG4HeG/rjKuY2RW3SEM+o0Bu2xQwtYOxCHuP6yPhS+OW04uKsv/1LPcs5yEXD4
KmogpTcLQj4n1S0CZCDZ3FmSez0GURBzoHQt2RU7UvsgE9uw0oTTm657BB8ltgnqOjO7W/TS3ssF
nYBRZWQ2S+SsH7PBsJOWVCIT5fUMcx0ABsq3oUAEXjv5oyY9H2oVRjCOGTuvOis6us94Iy/EHWm6
A8SIo5aQjpntuFMdQ+ld0CnLPEI3QTAI+6XBhTjoArvAob1vRU+CZ2U6eg8ji0TGw+1xq/khKWHj
vZCQtxYEXKRkNIga7bw7BGU1cCOOWM19zVf/wPg0QR9fbYhFuwaep4/IEWpFsrQtqxrv5hkRVnD+
8xwP1aB6ufquMcKAJc25uI4tpUJzKvn5XlKKF/BzWG7EYO62WFdN/06y3itt4GKP/eYPS4KJPiFi
vFWw/8/BpcCcvU+Q/I7hu4G0nDCBQBj0pWrymv0Y8rK9FePqPdl+ZSH9HUbs8k12xZWH+rWEYz7i
eeZiv6+hSH0rCbRs3sFsSJ4yGPfNb2sEKO9qVBV+5VvZ0cpikhmS4QYOUFfD5AcvcCkSz8eziCGS
kNPzmQJMzlsvG+4FZfLZofNTio2xiJEfxIcDiPPxrvk5+3XxngPEIBzW8tYN1FIwkthPEtxAkZro
FSIuus1kD25L00VoUwD8HKufP/+YeywIYLQFTMeQqQvlk+i7Hx106VkWylZzv2eUzb2hFOrY7vMV
xNtXoXmJeoznCSac6eL9UPIcGtg6DzI/d6D6iP3cUxMfRsx9NJORS7afTkP81oLihbE8z0t6MJTx
mA+u8IHR+o0v0eR24Zca7q5QeQcHmg4i/yP/VyN4AlbXl3xwwSeqRFlGqV2cGVLjOpEVzi1Bfc6P
DYv5VtTtNeOuz9eQXcmjngT3dMWRCQAjf1OqqQDzPsSz0XAQTrAbGtGkz0SO488sq/CTynHqvyjp
+zPBNOk2Wlt4LL5QJ2UYfL0D0HcB5W0qI1eBREh8I5n1skDe6wUTXM8EAL4WVzNsfxHi7uFvHbUE
4IaIj/BgmZuF1H0O9RUGT75cRk2fCVemjmwypiPimEKXZtKzVipfO4XMqaQERn/7roqkpGmD3UVT
+QId5M4tjqab0WZojszcMKSSlGk+Czc7AELIgFFAxkf2Nv1mWSTnvsrilGVhz1lZSP4aze49ylmV
6YbfSKqpzDcwKogGHvMVhdZX9fOYXtihMRXCqBVGtSp47AHStWnlxuO8haGdJygtG4+ZFYscu4Ly
gZJmx3f0T7SWt3b5OWB4UHSKq6mJYgYwTEDHMhymWtBqor0DJaLgHZ+Eig3tUVrCphr5lp/eUKzc
l5tCTXmafekwlohtGu5rYGg3PF8H1+4iNxtTapfL3Y3g0DFrEQm1KNRdi+Ka0fCH3duTnUIKtox2
go4sh57vEYxkJeis3+rCsv/W0eUnZzrYCN8LZlplZQSRusQmX/Equ+V6D8WXkK1RbDbUEz3EPQwm
lgfB8S5Htxnl3VzATgJsfJbeA4aQHSkhM37hJ4aFwrGsAaYW+CAYJjlsNKf/YfPPXE0UEC3iaYKd
LVKv73r1Wags/3zyptdUv0hfIfrMsLsA/YgwXSXDaSNbcpgG076vB/CBwzk6nOYa7uuLBOkSxy+J
gdrs/wGjqsgfN0MvGx0vamoHnnOMyv4zAU++EG/7TQuekkQlTutuTZI/1qRL5aFLc7jkQ5QRB2W4
PXUfEG5fXGh8CqqNAgtIVfUzGwuTh2B+xUgaxgFC9Ghr2rlstH3xNzv/yd16FWdpfUVFIYplVppn
6jCbG/OH1GTfAm10dL/Oz91CtkPoYUbiwXsZYYkkAb460HLFTWKFcTH+YLqrmMC58f7euVhC4bK0
tkuJQtTt/PjDe2+X3uaM0cqJRqhyc6KpaaRgLaZtW1OknD8lm/UV2ea5onoe3Jnofnjn/Q09f8DP
+SQTXGH/a1aAl4uZx1PQA+gLaE3V2kjtw0EEETsvHd/527bEVZU90EwPiBSvzn9qiu2+TG5TfUYU
V//T8RxJbDqi5lMWO/AKzx0I7xoJrJ8ZUkx00NdHOZ48r8AbVUUREOVDsJVaSheWsaTDQwp2vRfV
Wjzlj4j0yCBf6MHZ+7cEQTC6eflNGPqN7gY1DB6cJT4SsLLIunOeqK6/svJHPhOknryRqfMTxz7i
isASm6DTd8b7a/Rg/Zw1AgG79QUVjhuJCz37QTuIKYZNLa17GFbSAal9B4rv7z0r6bZChXY1lrn/
el5Dgk5j2OFTzmkAHL6JxHL8pr+w1ya/AlffRe0AHvWGgZuWo56AG1CKtyF0f4A1Ce/3te3oW4DH
8p7ounJahhDP5kqu1kQPatebHPo+kefPaLC5d6WV8mTtKmqbcYqYsifMB2uKPRjguYbYnjE7YAz+
1mZGJgDhVNHvTvwnv6aqAxgSCFdkiqvNeWZWE802q7vMGbOyHiUomXQ9zatII4juI7qVAZySVsas
G21WE3Wt3UzJUG+ebgOQ0OjA4OvMRg/J1YL2m0gU3RUXlDKugZYtKsYEux6XSo8w7C6iOmV7tGTW
fDSOqQVc6abSqPxVbWolaUTQdS/NG8EXKILCxs4+g0IOQZxfix971opuP2GRzwZV7cI9XJBmJXI7
k7iiyamA4AkoX1DIdvWDoFIzqvZdvIaWzWjxWcKLZanAmKyJ7UJxFclLkqqRdjuBCZYn1N7IoHdW
c6HNFbukNPpEqSWvmeYQoTn8ZaL66YeNviIJXWK9egAzaT4MdKhzKTmVML6PPaD2ixRCrFFViG82
zW5Myu65crWtGOV66fnbu5g2yvoX05hTd7kofafXN4TItOe7oahsfbcmUGicy+02W77zdkKVzXDD
9bDQNsm8jbTmVIeZ4Ti/DnARjEDCDM9Jg1ffdIoEncpQmKhTe51Tijhl5HItSGG8OMDvtCOkilm7
y4NiGqoq+s4M9T9iXoxqRgZsjX+45LdXVRAwTxFEDob64xZHHIYQSsPIt5hnKS5oEyBt2iW/UYXz
IKXucYgP6LOCiec8Qq3lDPA+LT1AUGWYzxclWp/epZXSmOUlX813nzCjZkAUggIdafEx1naOethW
hKY7ZcTNloIrZfgRbdqR4hwzcH5FZ5vHlYdTTgiXtbcOBp4eVpJmoR/wEtO8sauIfiul7zF24/cr
yUXHIma139hNntiZwfKjtXF+tD1dCwDP2h9UhsnRedGFcXlljVRKGLCZ4Dkt7nzbW7ZGqIKbszCn
3QNiJpSjdFHMx6kzKPe+iQwCuAEVssQibfriLii4LVTV7GlZxTIDmqhfcS3WxT1y3pUje8RDwjT2
6LR8VaH3E2lumEXw8kmAyBMEfMrmnJFtIgizE4g7DnDqAYB2CXrJ8W17u8QPDHUa4bQzNOQ6s9C9
5j5Bje3Hk4sQgPraiQ6JsDLm5bs6ha+vyQwkHaKL85pXBAL0cxpCoKsRNALoWzC0llrbIEChzhlR
VeBUdaziANeQPB9hl6V+ZGO6N2GkoxCUrs1ogjPhUGtM6lSjYi8V29hG9KRbD+QAIhXQkF/gb17v
yRRBfqqFJusgXrOedD46ZH/WETYveDYwAg7ijeU4jmA1SLnpvPtcLgsYb8DllAc/ZMG7goxpKiek
VaSNaApg/VvkYhw+uAt1Wbh0S+hVwK0TXvw2XJ/UAne+jPRvTZnBKD8NJQ4zZ48S6LF4F8g7qLoK
PKIodjKzxxfD+oPcDuBsFVz/8DOcTDDsM1w1/eulbu3Sq+yP29NHVF8OBA6p2LHp/0OQXmFkFPY5
pc2fAw6DpGymtZ7MkKnZcUnCnQ9ZMtbmiA9RKbVYtI/sYzYe4vaDgsjsEZi/Z9LSUEUkV9PB6woT
5RqItHLUgWqNiGJZAwLkEU1rbDJp2G4HrKkyfiHBDDT0Ew0Vk1Die0TkNiia0OWYw6DZjGfaOey9
McGx9KskQMuCPagb2jFF+wYO3z+H4v797XQqykENTYE7Rb1G6qpLE6xGnBX7GtnqmtEZ7t2Jilj9
yFoQUo3jFFDlNGdSCs9t6ej2RUg3/asFKSBM1eRD8ZAIc6VFskkfhZkgrH8FyBl8hpLAX9XoHgea
7fvW77M9bHagcVW/3OqlfmT0+nvhapVvbkLSRUaPJ/Pb4uVTdcBkoEkvZvEJ9KvUvOrGQQmiUTPI
BB/I6NvYEo4lTmpA2/dw5TOQUKKarKx19I3QpcSUGz5qKTGGoVvOjwPoujrHF01ZMys9EuoCUgLW
zKAkcQ59UJ0Ksi5RLFt0dZJdqZgfYd8V4tudMS7cfSS6HW3ziCnypabhhjvrorWTXK8OPVj97EMd
UXP9oPgx8+Ez1gyWHCVoUHOh78ExX483T+LRxZUxeifuZHHCViQ2tvUT1HWomwp5GN3vSDnEOCLW
0RrxMUXd8uLjigK+JlRJF8v7Nov4ux24lg0oj+cJaD9Uez0HBO7Lq5FGHC3bhzyL92KY0vh1qZLY
mn5xKTflO0Rouft+TCf1Se2jeaYT5nj1b1Gien3RpLwCsM/4Zc4Sb/VI2eZhqylSgrloFZzEh7mL
CnTpFV1cq5UR7hcD+AaplJ+q9PUR4PMBGPUM5gSfgzq4exOVjzVxwMngN06OvPmSUMroogUt0LxB
+FT8YTmZbFbLHi+aWR1xiun8eHbLOR3/B7H9FNwwuanebafIXnVRv6O6G3c6DX2YzYBYcnVG1Gp/
0by9b0T7GTL7miu6TOqMdC0hP3zFzwZ1Me9QgH0bnUf1HB9LoqU8FMZFWE+vXUACH6rsAkhZF2Yg
F+RDAw0ObvfmCcN0mxJ2Ymgwewsvo5pFZiXFwwlOyr17hgFPidqnMQytoHMqanrn29d7VYXbKA8C
Zd6X8jPFF5FIQitGao3LeAPe8NrTT8wu1RyAnD8/DBdzdwmWUL26N7qg2OosiJuI3VZwXRQvh+AN
QDnCZw+bHuDSO/i0LmZFGi5b4wxuyNOcdiqn3luLK0FJHY7IVUFE55r+Ac1K8l/a9W/hVxXfyc6y
8oDSv0AG8/Nl2bPrajOdbDPCDY77O4+hJReB+nPWDLaPYg2oPhJr8dWQtqeaHTG5bh8mR6wS8emB
XaDZeBzVEEtIf7QaavX1Sg6KeyrAaL3hu2LpTZy+YEOWfFIaA02Ke2pKkmGXvZLWicDfPMMcoljm
kSytiw6n5m/xShZ3rhckDnHu3uAa35CGZbFLGfb4eimEbkpgq7Jbb+Vkn94PBgeX2HFr3kD5BQbh
3prnXwlOkqvjqH9b+5VqrbWYUz4g9faQW5pMM8PwruKTKPcZ0UhJwtoCwDy1qu8TgTTwqEGGAS7o
uxIhaxpsdfn8M3G5OY7hxlBibMi/9p9CDtrn4SRJLVGBvAMu7rWcRY8N3wAwHMcRXgNH9LGGfl45
ppuxAwVKk3RFqu62VqIaXIXy1VVwHzpD5N8uwuL8f0SoXfXOK2bQwvU6HN+SAWwdRMUUowVIcP29
Ep2oMXSzxfzET3Z5I6hvQezcmhmx8EBQi824VaKgu7opAyvNAcOsu6MwVkOOE+yN6IeDMXhh6Jf8
CXQ0TCo/EquwJHn8xCy7bJuhstmn2evjzh4XQDM246EEhtPpyadvKBXChk0q2H6phfee8T2rSvZG
q5RClSObYt3VH3dPNkzjZK3AGlD4qnbZOawHgH/yUCiSa/QHjzHjfXmwgGmh9TXNKgvhe4tSfxHf
7IQWkm0HGk1R/Q7BuyIBtu3QtvqlEpQZMcaUvNHO0qqH4ehcAHFIQWNxDW6/IIfGyhqS7Hc7uv+d
PSKnzKkZqQY3WdAFvhqFiNvYwqZflC1SmePSIwAZpRJ8jssb+siYJk529imO71zRBeAHTUdYvcnR
0yRTjmKBE8hmfBDwx9/DowDvldlI/Ss4vVrNClFYTq6FfbyY0MBfkOdFPbUwWQ873zEm2dtCyZx4
LYvgG4yvgN3V+TnEYUsK2m5vgIWkX4RrtiKfUI2KiuXKwHxwOiw1//prWBbijAYFEFEbuHf2hugB
2w/O7a3J4jw0AGTMPD8CdyRqWr4lmnGMN3YS0TnQxU65UtHUYQtEEkxj4tCvO2/yfeG2u0wwicuB
kRCrBjK23De8aozZ5ujUio/B7OH/BIgrlUmUnOBTnsdf3r39fyP6bY5499A66GsJohFNUWgoRIkM
tbbg81M7UyKHKyZ8Rj27g4LEecTkdJivK9McTs/v+aszQgsf2i3/Q45yLdd3ChCvzyCcQCf6OV53
Ngb0YqOuDKFIZ8rglBtSwcCI/7rFCivp3INNEyF7BCuJlaJI0paFBLM9yODUeUuWBv48iidc4iWO
aSNPvCHIBQ7zbOU2JGNQyAOfplitA0N6gJS//QHgD23Wmrg0jpEXzEogOxdsWDaOWPyznBZkVIVC
hWT7ZZYab44neHwk9ttBwkRdRy1iQ2+1u2P2kg2SMf1FC3YqQgrw0ac/XabDlL+oi0W+QNoUElQO
j9Z6cAJHLJsdBuLwBOMFrpMdTQVTA41X1OgTSmWMIStZIvgBnNgzn9ClvRFkcSSOOx4/JGVSo0jN
mxtiSsuyE+opUhT0D+MpXi2WDrdYYK1OYRicsXYmBXkA/JPXdLy/IRIoAmx7/gUHajuGhdAK8KEy
Oocul1u6o98MBb6xnUDQRs309ZPF2VbMAfzJBqqH2hhh8/t+m1YYdOPodWt/v5MQSow0tcdw2gA1
XbwhW3xFHMOvgHLlh2n8mx4dSGDSvMzLFwDsEvuqJP9gy7vHkRXIZajnYR3hVcLl76AnyNN7bkRY
G7+SbeVhFjsWcrmArFad4A5Kr4aymHiyvEnqgrHzdZTNaG413nCq2iFpbZnsHwTa+3CdxDs6+2P5
PkRBdgWbZXVopmfdVXv7QP9jJ8KaGELZKvTdSyDnoGOumnS3g/zw71PZv5w9K372SELaIgwTrjEn
COFBYRQ1NsXZ8mFae6VVwfps5RqL/f1kNEz5qS/4CvLodOxqs25egGtJEQQLs1EeSoOhD99AEgbz
Rf0rn7+HawZwQDZHAXMu0twd2yMA30Obb6YSvtfZ3kqFY0A7+zVX2ZO5eqzGE2nFSButCzBiax3F
8BIhYpnSNcLpMKYG3fc3a85yLhj+3zEdLbgzd2mvj+zZ+yD6VxS0BiZk+CtNcPMjijKIiXW+BDhW
WRy9F1nZUmq84txvrXxXfb5ih3EQk3C1vHLCV662m/4uvKosdZU+YHAKVEvJnPuATfamy5MfMgHC
30TNb6rkQ3ApZSHfEyACtnXBAyCSo6f7yEnHraH/JeFEE6SaJH6roADV0xByN4pl4D/uTGhsJxzL
+P5XITXYVbf4VK6GiGuJIk/ClqkdWiItwatbZBpo0EoXH/BQtoAF27NmmhzyVWEEJxkGPO2m95NQ
iP+xVu28hl5Hn1z2C0E7xvVctR7M0aG8Hq/plhe5DXSJzW/5CPgf0+KQkD0N2xo9ETuEeDpDW9IX
paFhxYm22E6MFZeHn/bMmkv8EBnrozxGXcH5V5apBUCPbjITwqRQ+/RSvEIHK23nYM7qP6KEH6mc
3CSoneepJJ3IrwVNocw02bHSg3NIOFvdIPzBMX38+8oSeLb075z+IQ7XG3jAp5bCJK6/UWgGR3if
tR61LtxZHvdsr5qQ8eRHhjsvgq1pt2QiI0NAGg0lp2MpMWGKV5QZeWNM07j4hE1A3zaZbInWV7K/
71hFUY+GDQ9TAOVHdFH2TCDFcUVcdo91lGTf004W0PO1qA1WZEGGwNNCDFXDzHD6c0zNIkL6cTD5
idciRjPsioYWcgy12UBYPFRieEM0jxPm5Y+WKNcZHuODvV+3/HRdGYGjcUFdHMBAfah9XMM+rNk1
YnHgFExi5FN8+1yObqmLhZKHBEamzjK0/JBf7ffcPH1cZ9/v7p2D2pgkKYUfuwS2SfKzwle9PJSv
+vI/4QQFnb0dSfhXvxRSQ7XM7URO/d5ME/Obdi+izVzw+d+gHC9BbfT5atP5P2yWh0i5HcTiH3SU
Fg2xtMgYjKSdBtFcUR2V1N/SXTiQmfwUGlBlQpSojZCJi+YBSSmWasgt3RySL2G4fnG4PrcKJ2Zs
HMTgbtUYbp8WKd051swOvrOthfv9b2z2/8vgVH0KLxj4LYFqtyCvuqsGc/pK6Jh1C1sXBhDqXV+D
Iim7VO6cvGwr5Olr8kfN7bj51NZx9znlTtwg1b7AkJt66Py6pLQgnPG3VOFFjKmCYbLeE9LZ5okQ
jv9UgfwbHkyFna/TdMIgKayWtXUF+QNic91upctfUiAQrNDy0bI2KaZQIvY1/OsyJIFjjlAHFZ6U
aQem1ou+PcnuQoQjjaQqQZxM+Z4Mc+Roj2EWwu3OHZILjrVX1qrknkSp5JJZEKM5pdSMrmB9tc3B
TyidMgUnKGFmfgCUit9F7EACMJ8SIuUZly9BJV6dq7eqRiBCWzvTBBOF6EIICXME8y580YVzhB6c
+nkZMQLKjnE0qeuPghHeyEphwHjYckmhzU/XlwMYt0JnHYRE+MIAvfoAjT4Y0kkpVnI8Vhnvqt2n
BDx5o2bPuOUkHCbR0tkoCxxwaR2UiCD+x30zEqSQY2lKs2kQmQvx8VgU6qfL8MXy7agp9vMJsvxR
Q1NoBP61plmm0Zz2KPe3yT8D5bKWKl/U9nucNeNWOCGxlgNgaw6PmH8JfrYHTneSdwo13KydgQ+/
N0z5+P4+VEdTzlU7nje+UB0Zp8tln78XBEemsUfWp3OpFyAepQJD8dU7UlHh6lnjlUTl/m5UDImH
aeiFUkfFx3VR5XelXAC+EJe2SvMDEu7NQBq3hUgqL9j+QomRpJH4w6C488TFWmnLh4fj2O4BaJL0
PGLDa4gh7fHnI6+XIdSSUe4CxuIWb1LeCjcjCD7Yh1z3I1WP1T3VgjkuyIrllCjdx1aIiVpMt3Wi
cgxk4CGYPrChqFoziEvKmZsliocgWSugMdM3PiMsXPEhXJKdY3CSCd8g3aTEX+sxpwN+hb178EsS
0OHFWKxwAyDZZNa8kmVnUBxvfYUQf5/PVlj/lNvkEjn0zzqjh14EUNo3qCwHBhSgIBG+WG2evxKb
qdongJjnQweWN7PWiPCB2+EnasJLpaza4blFRd2sHy7BvaMGNiI9WNPVROTl26BvDwy0DwBU9MTv
3nkoJI/xzxm4wM4eKXlnjEeGOvqt+H/3FEPk/Ivk4l9+ER/u886Lwmko8KsT8w2YRS+/ZqXzLDfM
idN2ivDeHaqsJi6Lny4WE8uY5ICx/s8Pxue7z0uVRi+rlfAIRF7dSsPC1QAdQpv/RayWYr7wJ6EG
rIw8aM7hiOGebIv4aUKS3P+A2xwxWNhqNThI9W2dC/4g0qgDCVvCa3RcycAc+gFQO1/Ir+x0/9rJ
3Kz8AX5VD19NMFUstT2aHly8V3GphuyqHjVpHucTqKKCSEiUY40zXU0bMJBruleOB6nIM5+w4eyi
RoV1PBIXdBpflv0KtK7yf8cbBtXemgFmtpWINft5C3IgiiNPFbcQk3ISBhjvEf75NzGm8CUqYok8
jplWYl4MexP4AlrP4LjQVTcJd5IPh5I2cP1EhIA2lsdq0rIydFuTHTKkmW6jTzZRQ0uOKKX2Po5V
VPzbVZsKoUhhHH3TjIS+eSG+nQt8077bBnhmatJrErn/iKs7id+siXgHJTs2dYITjj2zakwuFMn5
V1Kv77eJ2X9Yq9zJGAMrZykoEPl5O0+/RTPObz98sQA/k9lYqwdePOpGPiHq4pCXhkvRu3leIfzU
KsGhK6fnWQWvpVhzFbIERnfcZIHFw93RUzseydjQZuP35q6ahg9udsUBY1Cg8pyxNARYgrvUbbim
dPqKZlqjvniB41boFbyJV3VckuovI47tvmmF1gdUlYkchUi8jmZ7a+vyP848EGBcyOwpGulPcDyN
+S+RkqSwVg8Ipg1zdmED+jJp9CGlC4m/YAa80jai7hQ5yZogahk1s+WGXWO3iAQZms7WMKrnoQui
S7dAicaMjBEvsuhrNpH+EgbhF7hWdYwZah6WXpLM6e3bLNTPcIopL5Is4vsXKHDX3t1qD2UAOoZu
u1FYhZ9JGSf7OJxpoB+TE5ZtBiBgwO23gwEZ4ztFqQkVsdjNCPl90XbtxVXGG3uwXFHdbAArAtnw
IuWarPuAQBMBaq1hLmqa5cH6tUBfxZuAKa3RASEsvOhVWdSYPImU+twSVwCOb/bLSGzlffasESDp
W6CWzA0ROIwPagiBQNJ4nlTUQiapumpHtrFn6KbfGgmr3mc6c95uo9fLrLmXCbnSEaA/Atj/W6HJ
edxqE6FXXazIoBW3intrSOJjK9HKu6ppZCTqJEFh9NT0AQ063sMQ5yPieS3DrtmA/165suEdvMTC
VDKmnFdeK4BbtJI8SFdCxrKhvouj2juN6fJ5ji1F7llKfVGfjASOO3r/GZ+HQm9QzUtlS2SQdDLQ
Xw4aZ18VLTa9iZhri/wVKVHkqZKJ73fZow0Ayru/QD3I+ZMo9eDHZS5vjr3s2HZ/bMkTjHRObACF
DfxOkNLSE5tVmVKsPnWWj6a890B6m8rcaVaZs643e+2LnoLy0FJKkVCClwy+UYx8ZiIELd+ZZjP6
ephheWiEE0QK1ecErhEQegvObhXx8AtmB8mWhMZj/RpmlxcIkJ6GUo4GxsRV5cr1x1hRiZCYN3Z1
ln6o6INkaQanP3cya+5UiLKpFFgYm6aMTBGoZAgIXS9uvKwMgpgeWNADc8fp5qLUOl91xXoUybcF
NzcA43W64ui6F2+PUTqlwo6XeSlF8UjRORduEYQCsXJAOImSbBw6dCEXnHhEPTDL+QSK5HT/61Fq
ZHQpNlsBbaB/EbkElZn9v5L8RHVFQmuvdtn+3Jz/maVWkPlHZHemeZPTJOb1Qpj2RFuFlx1i/HpH
rw851ntXHH/sTkoio50Rpc9CyRKUv36gSCEx9k6wT5eyzs5b1F8wsNqMLzt2jAaxnj19lIHZvG/U
MvvveqvqYBusdXzpKUa0kMZsPRXdyS0Tb80KF1Gcis6Dm2SizAAn0oFb5bMYNu36DtKd1jRJc08E
6TL9gCoeCqlCiOAHVL979EBxkKhsBlPGjUMvkQI/gqYO6yS7JIKOb45zfVkzET6apm4tIGYU7INQ
hruCHHSrLNvL5k1YU0hb9a0MUud04tqwwZB+rfLEosMgyPSvCLgpL0QLe0cQDP/5oD/d2+MQd4m4
1pwCsJJKw8fV8O+YHXdmp1lpgKgHKfB5rghJSM9yy4qbyGexFA57FQpyoOO+Pa2fZq9w/V5eOI4e
gAPI2AovijGtfG3X2KuGx1ypLOK79NcqJ8JT+SC6Osbb6H6U5DudCDJMUR3OPHSvQstGcCtdftu8
B01KhGlUrG0Frby18pAl0DmywMb/M/Xv+Ma/HnN74LV8CQ9OhrNouwlyV9Cd/vhMegNF86JbD9kh
/Sap/jPep8JCahgHc2pd9A10L03MyKzlrPKw7EBDAUPO9eATSJzxqGXhgHPLh4kNg1Ck3E2ye4vs
ciqlWLy7pq8ASrXRYSAlrBLvr4PVb/XwQb/lXkNjPRJCK3Yhwn/mstsYiMrxVpcCfqgwNoyTzSZN
fOVxTnfgAx5cSVyIrmG8Iby9XfntCfQW1xugyFv8lAN/FRMkjKgPwJQp/fhdXiwETrzC2iIM6lL5
sZJ+llb2jJlb3/dV0xTVw5a1DHyj6w0ilH9wfME6jrisREIt/CnNX3X3qV4izYZNhOhcwLaiu2qz
0C/yLoutwhs4jaEAk4ANNDHY3dGlLI4K2lhFvGEYF5suI24bstnUP03TiMIN2JNheWbsOplG95yT
x3T+77LQF3LuuMGWYlphH782rr+OP8vLo/RLLFX1G5HLM+6qnD2mr8YvUMBr2oVIWQzwQylb/kvT
dLDxLVUZWko+FYGOs8cVvgtJr1pieMPnyDSfWSmDSHNAflKD1bVYL55tjxuPZORtexh4/wLvIxln
HdblP//+fHxEOl4cKeM5NppcjNUB4BhHiGhBjw1WbqiWGsADE7TwOaGqaRt3GGtjLOkVawlVBonB
DDW8Fpkv+ITngFOFOZE3ZQ6QVCnAIKCkLIJKQZE3c3XKx5iIv8BM8DmqiKHDpbs6IvOCkwXI9a1p
nXw1emSSpTOhX9YtgG6cricWvnncyYlCde/tpBsBqeluF6hA6blybb+KBen7wJHt7jNmeM1i/ZKc
82C55dEQWsu1OEPFNVxBFuewlVW/uWU9xOKe/3J84A+O/Id13fev1CR1j9HGuoORNBZPXJJa3/cC
1fOyPopvnalTSqHHJ6bReLUJKdG0/3r3EcfbPT3w/4i0AudCAiC/EXIfsvDjLEuC+5PFvemsEpAA
Vw3QCy2sjttWuHgQOhOW9muq6+Vm4/ty2ZGIpRjtgDPoAfXpQ0QUycJ/S10QNLjVHDVvg65haVLO
mkqw0lMi2YUzMv5q1kMt6fmRj3g+tc+gsOYSr/GzJbpnmTWrZbep3j43j6fT0+2ubwn46pGhMVkd
BO6KI4tLE+UQUsHMet86kPbvFXNqVFyTZOTUkBpCdAcLs/uypBIxGuGkoPX9g58Qqw57AVdB17Vc
22aCrl6JT+q1pka7N8F9dLGXcOX40Dt8ESo5wR4aC7qtfU6GwEtZ68A+egnP5rDHOpj7XeesBQ9x
tnOv+xooesdQMlCUP5C6TmjAwS/tAmYGCPwMKv5pKCNljShgCtXjLp5nPiWNbshkJFzeHTs5pxNm
YQR7x8qJRBzpaYJzm/eeKutBqJ8ee1qHAB8tLYBgJekh88gYkWYT/uOIVNC/56yLlyeK1YKfk5Zh
KN1NsddTgVsxM+EspWbT8vJNrp+mng9f+60UV/Zq06OL8yH0zc3xFMnyiH6lW326nh40o9k66/zQ
4zRLwnGKjTc/B/ecYejFoqg73330tKL+BcUSJt1iFsZOlDVZSyQVrFLVu4vW3UQDwJIR5sKonf5C
IckZZgHM3yGAyn9ZLgsbK9RMkC846g0FysFKxuGBGlo8x0+tN6PYUhYyd/1Y2n1jcvJqlveN+RU5
Bp7mwtMim5+3yezmBsocA8ejBsBR9KTeAULcBBHyy/fa+s+uCdDAq6vQIMTfeO5lO+UF1mJ/Bf+Y
amn8+87Wdo8JYAinqKM7C5MWm5eLbr7g8kPIZML+Er33axl0rsXdDMExpTyLLbXWSJrLdh0UvKO5
TY5LUdlcUHasDFdMezIC8YK+0jLnU+bhleEycFrhqeUjfj4lnBMRnJ4/mbbY5LPRfQCBytD9kuJQ
Rha1EM4quiUvHD9qhDaOKVgRTWd3z+mdr2OU7a8u7AiNQjuALJLu3CUd154+CzcgXS5xL7FPjU+E
aB0HiNy0NZCwrtTaUi+lBAu3kc5+e6BRKuOcimbKg1Urg/+eu1PyXim93Tc73230q6TLLekvebrc
HiWXKI1Cmklm9c0abywTDlFASp0JXib13tXtuckZNZ+N/VWP4+7rzrCsghfX9KoGUYUWf74QrFqi
O2t6lhxj1AU4ReQE2e4U9vVFxxXFDPLdGchtQqp31v9xgguQqGOVrMAferZy4kS0RaYaLfyIbop8
OAvE3fH6Vw8VhD3yM0OIOVt7OVWDpY7S1oURgSPb32QKfxQxyvR2HyX0XwFwtJHfF0j5BNhg3Z1Z
7ZjqCs2GQXJ2nEzq11VPWHz7vbdahSQQFhIe0yvDIo1BBHuXoemtLT80leupTx575J5qnuvDaB9y
o8BoOKPaEYX72M7Z7vhD9WcQGl1L2I26wEhaHBbhGF2sn2WawSOmxo5OkGhtq3TY1z039sqfpLS0
kzvjfu/xhcCxh4bglSAER5Y67cUkLB1V1T8lBCRHChANZhVgHDd3SGiA8LeGYkSM5VAnOhU9SPA3
JUWHTE5DIrhYE7E+cNu/qHFtPJS7VJTdsxV2Clu8RcAR1f9MCzapquYl4sRC9ItvoXsT+7VUFPTe
GNLhBEq2b9UidktEJ1hnZUEK/eE/lh5hmDOneZ6xDtX+lG/7J/ailSf6NzIvKDyWFG7c9w0clkHB
Vnra/0hZ7dkshx/jhsbvPwXLNCguuqgWF9QoDFi809xNs0ubFBLj3fyeOA5sGbOhomG8iguSlnGe
8FmdrzWSflZ17KlqvUi6cTPBdI4ya/obv69MPo3bZ7M6+PahGJWmIzNCSi/tWDVG4Lq10qM8+KJb
aCOBSglWos9QJC/SwD6lCuyaWTyLi8Wrh3u7rCGxcehuayI5rahhh/RXfhTSOSQZVEd28LXf8j65
46JVGTlAJbvbKFkmdPczktsZ3dYVefCg/hU6ONb8eBmNQ7k9gmujSB1+ayxwY76Omw1S6Bxj6Fvu
ZarZa4yffBmyEGI8Y9jx8V9o44DvUjcljX96BJww5V5s95QF9wZ1HHuHcZf9oHiFH85744O+Va5U
T0wPEKgBkD+qQWgo0j2vav1KOCJgDn3qUHQUiPZXhstc7c7pCmbS7K5wTkiCAnpxkkrjydnJ21tA
UJRvE2hndtXD7nWLaJvJncjzgHSs0OUC+qgxRV6SkuHYbXMLeYziGv8P4J4I2isl/wppR+zyN3ez
i/4fmRupEBK+oRY77iIcjCInKkB5qqNswQn1LRnPWRz6Ige+5VtwK3z1vUXbWHT3VcgrKViZDMyd
b3ITIAspsoqOXDCTJpKLLsPMLUQF7IhLQ+tyWW1OgrnXyNlPx8ksaZ6gT2K+k2Zul8JOAJnw2Hn1
1IjChTiljbjuUJ7SMVtMi3e64WdFTraVg+H1Nvn3QarxtpzZrG2ecDSGgG28UoHZgxyyxcNXDMHY
McW3vtU1QGYY6OX27LcEvjmllLbf2yub/y40FEvIcd8AA/Zv6OlKTlFDZsyfLNL92ebdvhSeNU4R
VbWgA6wQZy+Yy5K3kEcqZhiREpmXMwquO3gI/WoNsxoZ9GfxMwz75i1zEU9eoXgsX6OpAynNRoXw
pL/J0JXvIkhUwQQeCOsKPJvLujbhbkUyb/j6OC07JEFqloQkoWv8zNAsV7CKzZ8gzkygsHPBseIM
puth+aaofHd+YQGeJL/jzMF/6zo4OJHp+3ksN/zdR18JZD327749oenK9t+WHLpuQ9nbg1RbB5Xl
16aHYfBW3y3K/JnFRU/pdIBn8J7LS/k2LcX+FRzGPn9mucxNM+zdP0okssHftjo3qb2YETcUybax
LF/K5KPt+PMzIyiwcLzp5WEHWWhWXkD3iMeFnfi5V83x+iFAULKhTIsQwp8CragKWoe0cOhPpUv/
jS7mb1qV9UKvBA/EN0f4m9Gu9Ua7rhTSU57ENULVKlh9cSLcAlQhnSaU4EkPaY/grLVvF6bKpMhU
lRs2JXsjv9y832yrP1DLPY+wdHFyC00B6vSk//I5jTYmGHgoGw7pGf3BmkP7lAECJBLzkI43xX5I
OOrwbeNLESBZsBllb39S9yoUiSMwCG6KXV6/RcYA+tOs6TZlc1Bn12Dia7mLKbTv/LXYCidm1es7
SfOpiUm2P0fZfucOXdzZ1NsvEYls8ySnMsRqvHk1RxBHqzLcxKTCfLQL9Fh01NprUYCe5kVAMFhj
AHYXhP0Gc3kz4HvaVmAVivmywVMDpYTRNbj7fCYIqOS3dVKTVlov3vUziqcxwracNkpCC0tE3LV1
m2sPt72rmSbDE/PBeqTzYTOWtJvA3efuNaixAKxHLXnxJIWmHftpLCO4ZS8zgh14CfgxvkNUfrQ+
xTuINFqe0jBwVW7oy1pcLzkYpk8NaB+TNxQrWUCZUMsdMfjP9AGeo6VeVRRlbwHmYfXc9t6id/Es
KPtz9MWelaMOX50OWWYnHLAJxsWxylS2PtrNWpVh22uDwpkV2odZ+ebRtbEodxjGekOYIZknEjKP
1mTg0PN438mfzUByP18tmZbi0hgbLpiuWLT8g7ZwoYm+QMRxdKnJvkBSBDn7ymKMZWoCR9dPzTY7
4m9zmkkq1UO79qjH+jXuNiZt8p5T8k63qagRY2epHwnyxR+z2b3e+Cdr+7QaMLVq5y8VjSIQ+Tsb
OjzJCL0Ba5+T7F1kC+y+iGaZj1CRL27SBoguhTk0zbbsMcUA4exCV58P3pqA1fqoEXOgAg/jlkGM
kfqYQz9WwFVGFK3xLD8BDVr+6rVp4klI6VUYhu7gxzI8kErwgyFBmVkNJkQBt70CNfSaJYUp7dng
g1SiEgwYilDOAzNH2mXmGkS44OCboAnZuqJdzVGwxKqf7bk3TD7mUDOmnZhsqZNaT8s2oXvHrW3T
XopDKQ35qPqkzF0s8TCLKbPedgZGFLyDibPObvKR49lU9tC54ENfGrIECUZ/0jMqeZEI1fovwqYP
Vd0UfVuLwbAgcVBDaGvbnHkSIgCyXmu8jYSo5Tr13tdpiNEVFo6Z9jHOYAuO/MJEHK2EOHtsT9zg
lZvSQnU65HNPLOxiEBoQNoBGN605l7kvMIA8tfAr+hfqPOGjMSMYeG7RYAGp172M7yGtZ3053dTM
CT086e93Gnok8EJKSeF46wLr5ugK+Ic+0djN4ZLc3srzEx2VVMsvlMDnLP0v2UKYyoiMdiMdKOuM
0oF5b/6xm8Cbn/yhOnkdaNDmtbMJfVmS47oUpqyHVrE56iIffblouV/qhTugHG0AUhs7VRvgS8+C
VZashzUkz9AQ0lc7zU+yIlSsImy2bLfr2HIemTFeqDHwRS4btudWe/vOLL4NLL9X8JWya24WR3Ci
p0fbmUbrvpFmuEn9phtccDJ2coqY9C4YA5jy8wuYZtpNCI1mugEwyfw1M0CYLXOVhnhesW6h+4N1
8fNtmylYkgPGwv1NQlqrfplo8PJqJUo1TPvFtdV8LwtGNVqKgtQOpa8pKIqVBm4VcVP0W233zJqJ
rYc1L86wRshV5Bk5kCbmHGViOdC140KKHlyR83qHzVF4qo34VhTyLl5t8yZeBk3szbM7291qwsgR
E7p07aIHweIrcHPTFJS7U94IHZ3dCtV6T51FJYd/u/XUE5BJrFnDPlOgT1ybpTY3EQ2eQ9WWlS+c
5x3RIzH1qk3SA5mTePIWYBoN7Y4K6JUt9SmdB/I3T5btHYjC6mcqDusOIpqSC893fFL/oXaBgbwc
88tN7ZiVUDVTu5ztWRpYt9Q5HpC+OfUoz2LHyaE5K555Yj8bwwkmSOv/2lWufdi5CgZfmHNHREsg
0tWi5aeDjDAgtJetrtueFwOk0UgwM7wtNRkMVmjSBaajbkxQxtQF5c0BAvHEdeGu09CimHWSjF7X
7vGnnvcufUDEFRC4Lik0wHFmJ4mif3uFHEInKNXPNQGAUi0R4RqXY0kxJj4Na76kek8/gZgdgxZr
N1H5Tm0HtPnCy4N5dUYUI2smnt6QeOhB+FT9H/9YbwXUw5JcAc+fkoxZwwClt7JKsKeiWBrju7j9
W6GckQQvFnrmJ8uvoouutXFeleP6flIgvDwpOW6p9gCKEhlJDGz/27szX88F5H7ozVGUk0jg4nsZ
sdwtAqSdBRKLHv9QPDlqn9XiM/CqxQg+f4G+qBcuIyWNnqDRvwWO6zV83uAg2CmbwjLswMxq18OT
Cprz9C2u665jU1yeb/yjzsHPQ7aGhB5grdGS1SgW+yYZQ2Hg6Rj3eKNmwIbq1ygSS5kA5qlLE3ez
/RoUtObSFfvUmpTCqn7TBk+KrBHIdsQc/kVKZg9kK+bCDuEniY+Tt6Ni13gfG72Dt+Eiw8P03bVy
D1fp2Dw5m870AWe21G6CUdwMtbZCL6w0+3hf6wOycBWT9FL1cZ8jPXt056n/nsGiIuGAXIgqNM4S
A4cfpj6Y0Dge/fxATIGb/MI4xC2NcTH4mTRI5AuGeWjXHA6LR3IjSIFJguGfGRt19dQ3MkMm4GQ7
2wi1oIjOPTyfBIiJAIHC/Hqu7H83GMxH66c0qECGbOKlzqgxr2EPf6NPYrQ9Vvvv5fBplVkFzM7Z
aiy/6YiC8uB7s+wxQDOZQl3AejrgCndDUoIYREYnSBtI8pWQ/C40Bo1u2VP8/x3FfIWicB3NnTMx
D3tAN2M93YQUN6cdJCK8NgxvEZRNwMXESYzJCrn5Tp7XEqcwdG/eY41iZMonYe7Vt7YNPoK0dDKD
hglIxJcGkmzoD4qgx0Dy4BHe9Bn1pYKLGeS5Wj1aKgxsOOlRg5XQz6tk91HVBlS2XOxDRe9ET0Rw
XMWqYhQCfeKOSthjrreJ21ROfpni1uJlXg3EgrGnEgcq1mSxJgnHWAQfVNvYLwi09+aWPf22i2Vj
lRuJG6syjP0ZrrwwueouQGx/Q7ftooaVWE5sU4RvdwehYZqhKrdLv9G4UVB2wYAWcwK9o9v5dUhI
cUs8sGdIyzMD3eJQSjsHTYWfiUxO2FDeklgjwMWLDMfjBubo75aQA6IruVkby7eXSQPKscicftX5
TLVlG6WGfYiOaK0ZttbckFcwfdqwEiNlc9PEI3S1ar+WudOw/vY7PfO4oe4mEZ5cR7MabO6N2esr
ynwflJfynZY2j+VdHYIkzHQWzgwwZbJt3/6SnVxo4hmwLfMtZFNV03tbxPxBhMQULRT9CQqgV6Ii
ElVj6ETnkyLauIm+ghxzoEpHVNkx+gZObUDartlVoul+r6LTQFAzYGE45rjG1V6lvsMqN8IdU0tM
JC1YINW1JItLaiVYpB6QWrxXD+Jjzgce8ZCfZXLwATWWNeAwXV7XWZn0ARegEvB+Ipc8XdZPjdu9
ghncyXqQd4iAdL8SxbHWhPVjGayckCjaHH3o9uDNtBebwPDMdk4UG3fh87sSReIrtM1/lkBCgN4F
GwYa/wNRNnj9VizVVqw4O/BTYIFBYXe5a97X0rWPqUBfJCkjeZu/i6SnGcKibC5LISxnc7HECTy+
FSrBPP8A2uuLwHActmBK1x9JEGtecywwxn+ovnaWOuWPHvmS+tW9iNJXbqsNEBx3KHhUDX/U+hb/
YZOHStjve3tYpUz29COpvfsJDP3URyj9W7bKvRsQgrQ8TNVkF0jimWt6hfT1dDMvxl5IVip0Vm+o
YXJ4S2P8estbA5p2saNaqJ3/4gT8sZsAZ/2p8jXBj9fLRWP1+WRfq0YrjM5XlCmXho2O+Ve7CON5
03kUGLrUI6SyzcfrLKtq6qj9AsQIRkLQeVzxvdoTBtuRArFa1KoCyIPBVt/CRiCwvFJCBIUSEM2W
28MPqUxwUFF8cgegfpC5EM46nNcSgVP2YzzNWtKi0bMglj8Th8Y93ItanyNbX4Q2WeW7BK8wStl9
H/g0vOPx/I11tjMjZ7iew5WXornjVPphR7tLqwY+C1hWN976yEpKJr/hco05gRaHH7CYnGt8Zvf4
mBb4Pj7t6MHlKTLtov9Oh8wsgXF6PEyESMCudwH3g2TOwSi8ljQpBhn6MJYQH8a1rEEERHmlHt6o
cwx/NhmBlszHy7skQIHIlrr6osClIYL1Y0Q2YyllstidBqXNnBAR+RT+J+z3FBOAzIGUW5LmyTYo
qLSyyddTC/G01NHkf6QmfjJq1jJG8grlFkrXm5eXNJJwVWqtnH8ZTmVSLAW6n3MT5e0MftrXc64W
KFkfoiTvmqWokpln5zd0g/3nCiIsC2wrYyfbQEJAggSgXSwQ0zKX2pDLdLXJlC/87ZO6jctu3DvU
S7nSVkuloCa8dq7hWzE05sYkvHMQtfvp1p94z7bu7NZyGDOnSeieEimq6lJ/Q0+o0WhX5aXbie3F
LLBE9y/Pm/UBCub4vHh+c77tReSrHrzNLctHXiOCl7tQ/AJVyD9AQWnBBCb8JceUdMhqDRvOytFA
Q+VgwljmiKNzCoizpyzjtueUbBFdUOuh4IUODqcb4/NRm+wcbGNf4JNhV82caN3+vEpQ8rz6elEK
T1EAkqDyHXFkMt+9H04w4UxsqW8Q/FLAZKBBU8KR97xnRR0QTCRZkucb99bnTO7gYeFsNkPIa2Pi
ZM2HQxVMpdQnZk6UhM991sLEhKtnsYOYuLFr7BBSsxOfTeiCbK/oCgvlImWIBUB7QPjaJxbvfTJh
SY8df1A82zhs2oQiwBlf0VX35/IvL/ro2s7r3j0Yi6i/bMmAuqd1pSoZOs3c3+P173+AzAY9mCIP
yv4Mupwm/PpZFAxzLEK86VBEvR78leZaYHsPwiE7M//I1vUjZohfvdQra+EM7nGxZ9wQTXKbe/vy
QczVIPPdOmA8JXft0kk8wt9RO3g4OZBH80yYMlVdYz9Im7rAF6EnWH8Wy0zJoSSokAqu5A5FffiQ
ZbEhKB7LG2sFph1C+pZlI0quYPGGadzRjQ8msplohi+0YYZrf0035nrGldyh25yC9nznPNYfygw7
piEVsF6ZChCVZwFzbN3QauxdzI6jK8nTXBiO2ohLeyq6GuANq06O1AfdK8CYROKOPgfrbnTJi6/4
FXGILN8JWEoxvJQFs8umz+rkfXBLbRjkIBEigxG5xKyDrYR0HDuUk21MA0PHhFWhlwzq+jCvUIde
+BeUIXm3Nfo6kkkOGpD65yiLTOw+QqJ5OBC9hSel4XroeC7aR3jcLf8Pmpkfn5GFkMpKJTrkX4Ve
TKYu9fLNaCln5hqRoN2F5/thYZvEwQ3waLk6zQn2tskJkknKW77iu4Or9CtNcQ56tjlfLD3b42fy
vErq9y+I4Ja3Lb3pHiSzCwXU1s1zxyL+N0+gfx/ELyuJSvDsluRtZ8zcz0ykPV2Fqsk6dWziKBDf
BnZCZjXfaVPPnj9X9e7/krH5mfVB3+nLcNcv3OWPtqO4ehSG3KS0yE6ZVUrom5MPLEFUDTdGXiL2
DCWoImz/yy2AaZ3TY6wESzDH+YzGrBrbQK+t/s1TBWjFk3uWIH/IDIYzxl6JSfX8iy4zno8aozS2
nLdQ4ZIQ3ovIx6E0IwTHuAyGgo496UcgoDS1PdbaUJRFc4b6hTmch6d2GGkKB9OxyqXR/YuLxHXg
68rUhgXRPMxSFrPjat9PSrXfMsUQuXqcQG29B83WD+514dCJkPVfhuMRj3tJ2AmZc95Cr/qLPr7o
ffNTSKFC4qnUH9OXz+H8WQf/Le084sAc5/KwAP2trjszlXJoO+ewAexM/s/u5ARgez1DEKpc70os
fKUSjXMZRAAN/CYY2VwmsiAhY8jC5p+Yuw5RGKM7wxN98psNP3lI2R7bJsdENZeTVEik0cCwBFfl
jZXnAbNQ+qy5fUbFUeAPO5xK51tLrGY+F4dMsFP/lN1eyUlsGOvGpo3AXUOlV2SpDI+rEnJm6nbz
Hm5COdO39edwAd52Sa94pRpEhvYUQCIZ2qFOmN7OiPs5lYz0d5g0L3DpsIc2nl5P05+BXecJXr6m
9L5u7Kv6cjhQ/V8c6MAe9TCRZohUAsCVDaWsC3+7ejPkmcsZTZBFuaQ522/+FrVZuds00vigf0Vy
FnbonFZA9CcZKsDkks7E0bhkKSn96LGPKpIW2SVrZsW3x7CI6ULpXVwZYC0cfK6vzuPlgWWc+68w
WZrJqsiVwoUkz75Xn9RCr34lJ41AQAjNv/qapCrgC+1YkvPelnifFbvyMRiDLCg2IBmz3JjEary4
gZlFDeuy9FH+WUBNwdoJxt+53Cn0d4lGIPFNOhFx27MmzdpUVdihLX2QsBs1ncnC4Sq/gxbiOXGb
bzrSuc9ptm2hfN6w0z2s1FuBIEcCvXSZ11ZNsECcayD6wcdQzU/wNPw18NZMOF7BVrVaoW5+oRvK
8AwYPjG7OTUGU7AtgWitOjXRKLN2qjkZTfrWQgbOHth4Ua3zjCOkKk329tZtJFvmohqDGzTvSZOP
xbTbwo5/3WFc02szHkZxJMbDnDI/EkExK9jZ45gET6mRT4/LjOKFUVFhRK2Dtraiyl5R0lzNFYaI
WjNIqJhjxBE/EjvmMRlaMNXKmaqbZbXKetQYXwAloEucNFIhusyl+yYbjvj6IQU80fQxZLdmKyzY
vIIi5cU6EszX7CjucCF+nF9wF8QgHVv7F8VJF+DeeqLwqxSCZin/ixutg0E24mmxXdvSCZ7Iy/5p
fXYX8tU3oM+QNxY2+UewWJLJQYJz7y4MFp2MFxuUmeyxX83Hp32eOn0oEl/pN7scNKZA+VC8rK/M
BOtTo4FHnIiPivai+d8xnb7MHBaM3m66G+6cLnwoSX533Ua8W3JPtJNqqi79rjK4lBzYp9kmYY1g
6iA2JnQsKYaf3DvWMgwBeUA1k7uom9PxAHdGzUPgWb4nwnExTZ4IgSTFbMz2a+2HfeEaux9CvxHa
wt+4khQvBn7xV2rmCGNfMkHwJsOXms3CGt7274mYmM/Z/FvUjhRXmFBHu6vRKai4dHdNt9wRx5LT
gXPYfYdbaCKYaQ8GTEd0hG6hmmjlkFqlQu3Pkopp+CZpohfpnU8ZFzBuCGsmwE+cZXBLnjAkCfd+
vCCzmpcEzkHj5MhoYNNp9BfKXQ+GuXzuZ4Q7ZInyiMDTd2l+XDL/4VlwYcwXkmpQ1QiqDjlvwpBB
/Xhs6V94regnjCtxJWyAyrr9W/QW8jFi2cfKZ3TQ9gLqzil2Mo7R20rCmArnbVXVhhimK7rV3tyl
yCqvVAmV7rDvE/Hp7g9pcIaRCGrB0fyu+2ke6JXO9wS1L/YZ36hn3PIWRClnOIMdDafs+r2RkWY6
PD79eS6q0lDPN+QQd3P2whcMjnREyjyCtFOKs0eDTuBH4BE3E5AGFexHdsKcKUJIHSdDpTNQmlrL
RlTrgQl/XkxcvQ9wpWM6dHP3sj6kRT5PXghrqtcydPCgHDXumi0DyPoGJnG9ZPfyjONZWLwrfF1C
PnU0UbnpZA5895hXH8NPd3lQdqYaabW5oDecS+h1mzP5LJ0khDXy7ud80CF+lRTLAhgbmE+Y+JM+
i5PQQeE8WnN2Y5WIcsWIuvjCONfjFB0tBbGssLmyWdbOrJi4NzhH6yM94y4FobXw142tRopXZAf+
GhDZORa/Chj0+7HZTFTNa/FbD5btg8dyWn+xfOAt7zgBYQwDQ6qC6Zkbw+3qkLtuyZn+IbcyTzHA
6vP8SFvYbXzciDR613TbkIbyih0TaDsPRu+tkjA9V1Pk9Ove1aBpqNFIuUsQMetIky2CdSpoBRrS
z7P3dfF/zA3Qw1TnqiBPYxgqL9OP5J4QUYd6mgM9HIyYv+5pXJHKkhhjcwovC8oPjzoZmuatI8DL
r61Lkgu6vKaePr4E3iUzGhm+5dJ4IIoV0V5XObt2HJK4n1O++B7RP+DdaNdqLTwThiIqz8CbESe3
H8Xa9SfjPZdn+mXgMRv7r1/64GUEJ+BqlNe4a3hyo8uEh7rXJTU7BImDcOY6xTmfRVzZlMVH542u
6wbEm2l3JiJMPqORnBEw2GCCkOOceHaLNIpRawzlyzfDTsYDesdqqWI8OFdWtWW8HJhEVQsyDCYy
jyNttrcQunONnMW43k9dPFYKptKcHfqDqLfusl0qmMdYc2OKpqdZwk/VWqIEISJ0yoCC38lrYPJb
qgpEwpsUzPlCjoQwxIuroIPga4rLl979QEOKEadBfDvKqGprtj7E3NQtUjtDR0/4caIW66a02woM
dxaCk8rIUp4AbanJgJC3BWsaveY5qejQXLK8VJdW/kYWXQxoyT/jFYcCMsnLL+nZpR+aNYbyOsac
sF/W3wOqrzuP17jRfWfKiG3CGYezdsAAgAApwQXUIrgKc1iwf9dLPU88l7LYceiPBDK4gWJLqRWz
GsAThFMpQO3M2g6wRc4hoZEqp95O2k/L/5p0+MUXDyGPyG+Dk8b0+I6iUVLZN2sDCd1IOlh2Jw95
ozUwj4LxGdIqVv3RHNRsByVnsOQV+WUAwyAo6dQLSPkUjIstutfhBTZ/g6nyBKgdYr08mrfQw346
nIqgD4NmTWx81ilHOcBqA7zSzFE66vqLKHZ0Bt9hALUJjYNNu6tQFwNsxQGQJsiww8q5PycYsGet
C6fztLeQLvGqEMnIhbWpK38CLU9ZJEZYlJBrQYbpn86TOY1pOXaJ6UwzdYdVVdVWAtgdpXx/Jp3H
G2qhHmiR6plw/eJ6PpmYMgtZkHtP3GDLLoINYB19OSxl7q0UGSLzVr+wF05KZiNWhOV69T6xB42W
DGwxo/kvR4OK8NGlQra7qb9ZEQY7/4pwlve9n+dtlD9wO2tvYRyGhtui9N+BbB8Y6b6INuEOJ6yJ
AktAY3urAEjSr1r1a62FKo8Ycr4C469SnL6AeXkKSLmGumfBh4Ad2PUXTUom4/4Euk+6ZCiZyjwF
RcDdMxXcD5BgGlaPPLF8i2pwReT8JQlYTbU7//kdpNiTeq5E5qlzEEihD8+3tNN/ZnIZSVcGQqi2
9vKk9ibViQ0LetFQi1NZe0vL9WtDOD1qO+LITiHY09WfJxpYxwzsPYphiSgN9vSXHvVyDbQDWwj7
rpYWTSNlaDEP52NkpJJwZ/Ddh+KCYhNwK86dRlux1VCAi6sr+d3ztMV/+qE6t56kn9ANS/w4oiSM
VdW1CQhBUxHI60qVITwRP45QXfW5FuOYq6NRKPLKiId+t4psukLn8TdWEySLXYi/KanzROpz3oa9
xzQH2toM16hZmgt2VzmLNq4N6ggIAxEGcIje0wECMSqjPZAKPfvHWYWUXU1JORbeiEUmmByIQaya
i57fOs6utUBhpAp4RnF/th2KP4k0jiyS+r2juQUprRaJMnRasbLGYz6DCD+6YQu8wt+4HzvkPDMv
IuBhqk0zeF3mlvoF7JamZRtp2uC8uXomnBmciU9BhTiLEQ4g73V9qVOt9wU9FKcDk9H2Td3ke1gI
WfXksXNEaFbflUPoesk42iMbpdB9jMKwyPh6YjFFonEZZjSLrKH+6KRqUddzsTDMnSn0y91oWlxp
spHYThqEUxl5S3uh8E7+zQVsZhnNQjzD+xGvFy1NEP3XgoCs7kaGWoM+Ux/I9CAVJjFdoOYq3g/j
WNQe/h+5AN4MX+4mJumrGmtpSHJVZddUa6YOXyCw1lcs1vHGXvJqdxWit9RzmhEYNuiFPvKUNhcf
uVFFC31H5FF8Nnk6hR3AKBf+9DuisNy2X1tkC66TOJ4CVFTtf8oUxsZCjDKu8ymrRQ/WmpbEQEmc
S7WpgV9zxPVfiAe0yBl3PuuH/P8R7nOpNaRr5MgRX0zfR23vuRSVqYsNywE/o6i8NMfML4zu1SI/
NNqkY5+IsQTXZJZV8mDxgQo40ZZneEKk2sDkpScyj+5GGofSrjMI2auvYkp4jVsWoAlXH46SgvSe
Ae6MLx/MRbNUhyxe71CbKIBG3IAjlnwrQTZ2TKkolS3QmQ9vOVGUmh5nKY6k5Qf2T32zB7uWPz5+
vOpy2FWsMdr1VoHoLKtKALZZFeEUHPpsuk/h4sfCrqS5rkB4ksGcBzPJP/3TtmulDDSZGzAmz48L
WFIp8r+OS9/6j43WuZjIPDGvMvwvdEsWijuhQ24VPJwWWleUB99INhOLXxeSvlD+TEmoU5Z9kWr8
PFz853f+udPaHERsqu2Mp48pN3PMLiItiY25Owy7QSdMRBJeWx9mlVZHlJZqXjB4MelMk6/jeO2m
PHKY/oSZnsdXMCj9G6hX3VPRaAYKVIB3pmIfnrlWJS126zTIIYDuSfeHMxgDh3Dzj8hM79qp+hbw
furYZhDNqBZThgDq5srj0YXGAJ+qpyDJbkCOdlEPCjW3+8Hfth3c+7poof80QXr2ZFm8HgWH6Cs+
X1HnnTTRkVXeuxeuIA2dxCpNwrvTtTp1P8sAcsGcYl7Ybn5l5fC37pSJYqC6UKgG9pBe1xwkF417
mV3K8yMK4YqwlQRAaspfFv/3EbQGztwLv0Dy5hejKHQoSSzfIo+oYfL9Kw8T1Orn6TFu2ItLRiwQ
f8X8tI6l9WwyOJeTZnTL3h68Uoc5Tz0kfEoHjAG2AHQ8n+wfcEE0dwdIMob8pYNwZP3SjhnCf0ey
ypHYzLfSRXAAquiJXohOHWstBayW/nk7tnPdWsq/q1QzjZKdsJNUerc110KNV5+Zg6YE0HK66u5b
/PTrzgnhZjcm8Zk3tJtbknq1pj017o1UiQGxB8JAZUe2sOabmTwd8lVzMT3qQyAlPOPwFC7CePu7
3MTXzW2sBSD6WEDN3/XjxVGYsCUREO9SgJQZ2q0BK9AH+EbjQid2FgOKiwYAEGoa7RMVWwGWZpaX
UAE6kfwLwjiXs2Xm3I0rxBrZNQTO/dlq64HXmFSiq1dhC8PLET1h0P5cVIaoQBLqNTnTy/r+dQN0
hwzohP0bM3qJIBWP60yXY/G+vGasghuIpY46M5GZ/iYsjkiHE5xHoIbgobdpd0L7lBXsILZ60UDP
fvZgW8AhydXwxypa9ABpu+RUg8y3QfcWP1gFkjA9cb3sljREWTJGRyyoJKc7TDqnblabIZdvqj+s
H0AC3C8zw2+MNpY40smyzhz6TaOPRQo1gtmbjytnJnrSmbJSwIUC/rct9ysbuZjaOU0f/+8OMyD5
WUec+afmSmyDVvsF8hCOoTudiDKSrs3IZortKz3ThAcwjMdEIsZzPHW0W0CqZtrT+FoSFymaA9lB
eGJzdHO732Rwqw2WFQUYfFA17XRUWF+UOkGCNfir44UgyevGzfikuGi+wDyKcm8ctOMNf8Eww9l+
pmlquLqNdUVvjyhOHXsUflGNF+aoerBKxVu53jn5sFvrpiG3nof9Rfm2YpxJABBCP4t+h4mobNQs
0Lbbj5mjD9cVvWOKENv1nYSqOwaTjbmiyNG4oUhCzu0Jwn6nSAYaXjMBdvQcwedkjpFiLJy3bWi9
odaPegZbHQJq/MqAcsHzQMjDq+jJGmKEWWl2yJQL8VOSUdUKKn9irSD7grE66tcoOn1wY1gbNJJE
koZdCEBXPeVwdLucYtqFGjLmrhLLTniNUAHjWkGg7uw7g6yKsts8aTAVGQO7of8nE7s5URg+fuoL
9phcAgJUYVj8e4eaSmnTb6r37M+WtVq+s6ZJFTEqNrrwi4XmCPiokYF2D98FzUdqZOATwQ1JzWq8
djxIYSAc+ou5LSIpmtg07Lq/tj8i0d2qPmpEM4e6k/kF/OukzKj0jz8N5fCxwgqsXLC3HGDZC3F5
6eEzjmlcr/EDz5lvt6zgrmGnC8r8MVrRkmcUUbEoafRpu2fvMXQCT+ynLHUn3cD9dGuaUwTKDPYo
TRdqzu9to5Hu8QFU1WqJcQDN5K3iONqrBUHb9PZ0rQqFcT67CSqAZMh3gJjXTc/2dkMpikacCJIl
S/Ylmudt4bmzPaNhh+hatOq70JOKS/dKHKNIq6pUDco5hXuPXpuy58NmNh+rdDJZpzJsj1IYCtDk
M22yGk77xqIzxSVlUgOmiyTElvJEPTpArVwOWLOmAV9yLgZ55D4ZGp5CG6RQFoYuaW12tEcczqn4
AegSry9f6/M4GStmuZ0kCKJVt/Gr7L3G9UkEPtRDl0rhlWgc+kz5DYOBp8hJjfmOrYokEBThJrHK
9EUzqC4gXCIBDi6Jad5Qrf0XzQ4kAyxIRYm3TotCnA4nyjbLienvCuxL4BsgeFrPMJKOyc/tolTS
DB/ulhhS/F2+BkDYRNTVHLbYyYv2UMb9d1L/QqGx8sAVGH6YXnnuXqsa816IjWskf+6IEMuCbPxN
7mXUzJcoDqzuUlSv8lYh1qgFcEmZHIWfebk/HbH5VWsGIxWVRoK5GdWxvMIvhktqfC42hyEh5lz1
gYfLoKBH6SkI2kE+8cZyodJ2pzoWTPnHvAfXS22uIG4qyVDjyoCea0lznePg17A+DY8AIUGVrP3A
Wb6qShSOMuYQTlKmWY2y9DHeX4lsYETfc6eaj9MIRyvLwEmDPjqJXd50lTIUYUHzLbGAZTN+IsIX
me68e3oLJxNJJnetu0o8OOQ4juytUQxnqjaxLc58Xdq/TdShwr5vlvic2C400HfkpWdSYHJR4MFV
RgxqIRiI1N+X++d+p5JtBSQwTrURKVn/ja/7UM1KkvgpEVT7pUsWqRtk+QdUnqJ5S2CQt6KA1Cw5
73MmL9qbyM31Ihkto6B4r6Vrjj9IM/k1D5KL/lUHra9fti2EGxjQjPMleI0LCbgkbaG6nnLRBWLk
EaPiq4/3ToxvYiqiS2k5czoYtfGvg0aZdP7f0SplOHKBdD56FRa6c0u/Ty7JvawzVp5rYMjekmMh
XaXNnRsF2mm6xvKyxrSGEWEgtX/RJ20mQ9HRtVdt9TNb3H+c2Av8uB3SrZEERXV1f0EN1odQis/a
7C8qG+YSfXkges9WnD+DYoLWJvVusAXTD9fW5hXhE6IOD07yC3WRxjbaQu3/7icNlhfVnOvxGlwz
diGfDbhHqCUlEtNrgtr1HLgN5vRSmxi2myeLwMsgRv45KKEjCEYtubWbuIh5Hl+3rgEYIrdAFJX7
x6LPDmRbmeTIZSl8JeuqA6qxncezcoeTpxWJ1YAJMkqfNj5EIgu5+jLl4c8+hD76rebyw1YKkcXW
wgoWJSj4gR+7eyNlJEBAJvXkD/dH0C072jJYU9A91aTycmcioHf0pdktfPAwJoMIT1qVRyHT3Qal
3dFI+t4JQuxTRkI92pmL7v1EkLQQeVSWmY75zomhB4jpQXsssaT8cJEnCHdWwKtoECJakF2QDcva
VwB3O/6MhA2AqCzzbWu4yBshxSX6MNPjSysox12SP3T77WgzdyJoybp7QLe4YJusa+x0OhLkluod
jV7038QdzhU5DntWAciadeyiFIrLqElOW1+cRVF9wvnjEmGWi6aTOTOgMZrmk7qTS/80RqN8yysC
Y2QZhuqmGk6BNxPeZjsb2jsgAtiXX4hBnQdpe6K39Y0XCv8/TgVCP99+2NyyoyWNAkZ2MVDaL52g
a6OpzsyqsxezH+4zbJoZ8wQmawL4Q25AC1/Ykbnb5fo9Czg5SG9ipi3ZAvngmVY5UMNq9TcxsubR
HgtCzQUOrInJvVFAk1MKY/a9C66hVirr8yZlA8+DKt1ryxRdEzJmKp4wwNz8c+LPBJSLNkBqdoXV
3hkQk8I++qmg1AYfpZWS9kM0pLzUw3YTbnAjzK2hUd7VdgJ6FSgvVjbE/DiogxQ+TzOu+678bZvM
FZOllUU0qiFij/rqkJtRuW1VI7vtDLvS0o4ulw506PccE3FRuqBK+QGfFwVhjP7MxJa2M3xbtPgS
lXEoQOUIO49Yc2dmDDWe27CwY+KjbXupTz/0jjENbwGYDhFKg/Q8S+vmHD85RJBTpSHCzC1/+jFC
Wyv+HeqlJm9IANdhQoWNC09zFgC7treXQFXcH3H/ou7dr0h0H+I2va8U0V56OEgF7jZzMKGtXK11
+wffA6Kcp0NxXaUI0wKwYMV/8xgy/ZLW/qlWe1X/QCychHONkcp4J5OCyUTYX8RhBoXI8r+XcRYt
qxlDHb2hEzzvgzllD5QNDMffH/mpeGGqJCk9yM5IK/2BnaA1ttb2IOFTzcL6h3QZsL4e8OLc1tX5
SBVdJha8wz1WdAA6xZe3Vf+Mn2gUuW4fkCNScwSTf88e8T3Za928QrjqSliQ6VKRJ1SnOzN3VLjx
OauVg/h91+Mm7TaSg9u4IoccybmgqOOlcuSejH58qriSYs2mTxKlpeO3U8hO0OvcAwLRmykgcrwh
d/iUlcuoUx3ZArsDCYXhbe74o3huFGFu9GJLEMYLWJjdDhKiXmLYuegapOAD205rRKFNi12bPZr2
L430+ydpnrp3v+ohcLatr2nTrI7w9d3yGssNIpstbL82kzxS1DQVjExGuHapJS8V5t6YRCEbPu8D
pSkdLqtSDCQ6Xbg54cob5+xxJICdhYrK/Ru3q+dPg9tovqcaDvb1yV2fMwuTtE2TEGRGITdEUz/R
7+CLO6IIj4B1miHeRkFazqKQdjEeeMjJmES8mqaRNd4eRS4SqjCd6X5iWX6pfTEYe8ZzU1430G5e
JPYgTWaGOKMHtK3nFVzV65DXU6ZQPsThonJPztQLu+sELemKh2aZPKUlz64sRIQUe9AskTCOFJlk
h0OXwd/ybJjsPGm+ZvCoBQuL40AWLPmVZfIll8uPp01iZzwry/2qwPgGOEhJ/MmCsXhvRLrQtmmg
gfvNi/Cw0WB/auGaa9mBzdmg9KVhr36EDgHmdo3cr2imuuznQGbnZZKWpHvKPo1XEOTFCV+/Drx0
HmQAEBF6Ppn6BQCCn2HEK/9QoGSiq6RnXE5nb41M4hh7fSOQRiIU59pDb44hrN/jQG0K6rQ/+R88
USTpXT2USaYAgcRy20GbDhWF9MqPxWguawTvxRy6SdG9mNJ5TwTmXbJ+nE3k59UuQ9H68EdqCkYv
XHphnzFo+MsDzGZ+9biVmpZN3/TmKd3W517g2xOMd8+rdmiIXm4jbXnbmnSbf9KqCFCfu8+na8fv
cjIeOiC1PNqxOkV5u5JxAbx1ivLt54GdIKYZcfQsWBUbLemWZb0+CylC8zAaNDexpomJNR2SXj76
GmJ648xwrrVENjHsmSb/hGpZ4ENx7b9b5JMHRungRej2i4Iv5bQkr8q1KDHuh29UL0LH/Hu7Rt2e
cQatJ2BPDTSj8jDFS3kr+XYkGks/9V0VMgw84Y27eU1/Zv8eD07k92SbzQK5IxLxnacYg6Z75rvm
eAbZFn7P5xToaVyDoW5nvVFErG8xlY3q3Fqq8PSsqN8RjfB99wPneYl4AnSLPdCydS4ibCuseGpZ
afmMEA0HyH5XMVDO9QMhFwAcI6m0YH2DvziYLQTytLM9ntyACKlwLeZCKDN59tCF29b5VlVPZeLp
ZnYqjHEUFUsvNuQslRuuxsDpvEFrNTm+7wbd6LMkBt/uHdO1Wh5rSE32pD2Rjia0Eey2YBmxupAZ
68TBEQN3C4iHMTp2ZDxo7MSR0VI7cXIGkpnpoWeQZRQv/6p7ChLRTnqxiNZ4E07+TaojqvoZ5B59
V9fYjszgV5QynJZm7qXKIbzJxUnnp/nib2WtdT2yC1pWL0jS0Ux/xRts3aLI/MgLOPpRGpGvoVYi
bsdySkuNJEOXF201kq5lVQYRpk1NAUmI9roE9V2+qpI8bgOxxmuucuOkVEleiud3766CEx4RAD7T
m1zP4fADBkzUvPPV+IATZA7A0QcLL6ERNvWkW7e4kV5Oi80wxPVR47PUkHY+tYxGVWi0pFuOD5mN
PC2Rez6RUx09ASSKdtFXFw6OovAt08wK863lWhfFMX1wdHO6IXEvDju3DBIyO/HlpuUX7kuxEvKt
nDb4RUto7gZ5tNgEBJBUVg6K+7bNW7QHsDqwn2zNWLGXtxa7YAtWqdXgIsIFleWKQX1yDtHlRdIk
RP9mspOc6Xi5WVq11zlPyGMuGuMAMMl5fwiIqdm7dT4MpLm5Wl7/IQKrGqb3KwJjtbhPSVKPKZg1
BhEqx2KVoOff/nROnHIibftj0W1VZiwgCuLdFMdykB/5ZL0chF3W2LoVwypQgg18/Ad3nV4YvcYR
HRmRlU8oik4ArRAGfYjjhH7khsgFH4yqBKOYedbRUp00x75++cd6ajbWInNgPKeyy+tDln1RMn4u
qlrCAhuZiL2zYjfaC9Ym+3dvq5g9XMAkPdQkljviE0xSzz45NpyvAGfZ4veIbFQBNUGO+Wf4iMdg
m+YRqsWuJlSLnq+QjYW9NCrKDDQTMBuhV8zJxVQI6bZE2ZzaeIT3JaMXRbe2ks4OvSmrYOuU+xdu
RKJt1f8L8xHT/JmkLFLVAGk0IICeHtzjZjX9T+oeAIlifJWpKtgpiSj50aDO783DE9zc7aX9redk
0+JbP49fFP7Fo8s6bLSCmI3YnHzePcT1xeSgc/Ivo3h/dsa73xxKF6JyCv7801jOyf+ibyZzVwTV
3rD5x6JRu5bBN1iNvFrbfRMUzfs44Otwxb2e9oDvp7nNChmKmBWxNZPZhyIhXi87vUYudF3jWuKk
bXz1gBPwqf9uIhjMHGGnrZDMFZ3d7quoXF7ZhjDnnClRpZ+jK1J0ZT/hYyOBrqgpQzphDSfteyT5
WjiY2KMXC0W478d/03uDasOy7t2xYVfDS7YDNBCvGhXhKg8UEYgp7mwqg2jxJ7tYreM6UqbHAqLH
hyGL9qqybzGeVuJFL1bv9DRUQr+5OcUsF8b9Uu2PIl/1TJcUT1Stvf6jY3FCUehwMS/jWLz6y3BU
KBbZ3rIgGmIuP6jhNF9I31EStl0k2pwnpDDgm13fAxBE4hTyYnk+eUpPse0BR667lZPCOhgdX3+L
LynE+W46/e4jekmcYuU2j3iw+89UJhiTxJ2x4h0Sle6NVucGZIwd2yNHYb7mxsXX8GLC+NfXlX2d
ytjkkWASznN1onZ6TYA+7dScYzeiVrLMGIboyFOSSGs8SVG0GdJrvv7G/TxDByA/KTIp42/z0Rzi
0jOvoDN7XQQZYD7RvIO+rANE5lze+6d/SACCmaZhgsNVftsajQcaR9jhbHw11grvM5tcDWZ6dtoq
MIV4eNnpERZymbHdH8H8j5b8PCf1Fp1LsM48Rk5VNsbnWvK26uZuK9o3Tv43CvQsVcz+nFg58fgC
jAtQ1GA2Cq39iweT/cUnJjQcumiZs/B34p34x7fvzxVUcgF3+s2+SM1T8GJIoZmonoVlEHQwh0sN
P3SG4PkH9qyuHOwvXKuZhQAjb6ymerQylH/l11DIlYyvKiqhxgYEAfkUXxB/XM50OTwmz9lxRIaD
S4sMCcpYevUHsVEaHN8wr9T1WywrkSs1dm92VlnCBdMIQKZTZdvDyPbzOrmU3dg2rlry93NC6yTZ
d9/0T9wkBOyG/iKfdXok5vZ7VnaYMLVTy55RVH+lvTDmnNpDQ8PePwPAqW8xzNrnHLbyhlKQw+52
frfDkQVX+anbontx/GWgkDkBTedhp/isznXXlk1zFOYfpIwbNbsyHGqT2p9rymMgw1zhFC9w0VcH
ocOO2qpro68+HILSSV4+De8m1uoxKVRc56UGxYtI2we9gJf5MTtViE9nzrdQZzaZ7+k4pykIm8/Z
apjRIFTQaIejraLzttAH0W9x/4767nyyPrqpy3oSdRDzbzfLhNch6jJl89pERdPPEtNomRa0xO0d
w/9c8kD0180DjkfmXXf3+HJYhNBjlfnVyxYSHbZv79q6XDQ24eM4XfxS+vyG+s/Dyp0a+X/F+1tg
fhUO70FYK38HD8krW8H/BUfIynUhedCgk7inAj3v1OO/6AxZ/CIm+6/tyaYVSI3S204CoFzIVLsS
LhHEZCaNdE+JSfnd7CuTpfsahun06uQTI7t7V6sVMvWBgq6CKk//75FN9yEYuiT0SHJ37TRxwBNJ
FU4yo1Ry5uscyN8IX/KyxG6Yjnh5S583BQqNiT+CfxEzT1xBVjtWOHm84tU/VTDcoqj6TfQiWR/0
EuJAx6xskCm7Q3guhKr6x6AldKntvPN9toeX6Ar2QAM2HHHC4ZU+vaXhoWcMv3fX7Xb2jbObkiVa
zy9Ti5S45qCkymyOttBSwkyLN/i3nv5+Snw+6o3O784Gy6Nv5K8leSNx4XHjnh/XPBSbhqywA7XI
enj1Dz/XcVPfVjZ/8EdGDLkSUi33HB8OeWFAKCJEDuKXYOO8Zyj9xbSeuL5jYTH3rHdze9INh5/4
wCefEylSINTEWpKkAOcUSlAIF1ttzDUKv+YdwMhkGSIRg2M/S5TIdfjPiHFIacbSMouGgB3TywGe
vxrVDz/4peqigqwbQMKI46YX/tni5K4S8SBES3DzdQq73y1GEHBG0YwBrywdwY9DcZ71ZyvtDell
vN03sItl+z6F8ij8Qhe+v63ci66IjF9luS2CwDQenbmPN88tchRVEbswoMxfYbkYqifmZFOF7Oo6
UsAfQZj+4tFuhDTe93pXVK60UydfAYMBZB/ZTGIi1WwC7djaziMULet8vrKj4CPUJqc2l05CNGgM
X3WOdaU7qs6FoCeUparU+xG4BodDI4NACzsVO5z+tZYGYhLsLY00Njlkwc3CoHTlXzfWrcNXKa7Q
rYEXCJWKIDuk5Pn6hKHcgErbZOy4Es97lzk+3BsbCr72dt8ibbQ+oRVX+g2bg0uAAb645RwAEOV9
G5zb+e6Of1YEOuH3GDUg5w2cnBcLN6/VjuhwwxU2OHAkbFh+DoWp9mxvwwEeUXGCXf12V9H0j23p
JHxHL3+rkMiSuv0cGQHvuezSKGN3GIcnC325H+L6UFQFWpmqX9JXlbgHqst7KYubztSkOZhFO9cL
bV6OKpObXVdJg09RzoI+oImpLka23WJ73YeL27RbbCm9hUUwgltTXhTO/2AZ1yPhDPF1ccKQ8AYb
5hQ05SUCk+KmYCCx1Hp5QRikyA6r1iCwZ5g7YDrkcobpA0Qn+4Me2YDjF/YjItUv/75FaYfQOHen
2j/2ZclbrdL66qNpP96W167UMria8/NkAIXZq/Pzs4CnPWWFAhr6Xrwe42EvnNIgEIinmdUM8a2+
AfD0NMHFHHQ6XNprqIYMbKohBDO8ae9XXIrzA1obNxmLsQwTuiQEpV8+vUGGJLjvKkxKxOfUIhHd
kGgre+80vw0uPjYM/HSsh69zlduSMu2HuJrN8Vym1siRnW8/cp5SL4W0CvuxId7N5E1knpHn8sLZ
PFIWcGEv6VgmQsRvzH7bxq31uclOKQ8Ojck4uu793klEuZxJfMfuAYAKHPRMUjq36v+Og6KLCgK9
OcOBbbUQyCQv4ZxsRA5VeFbTQykT/1t94RfRiDapARBcbrw+01fbwRUl4xUDwsjUBN+rBmNBHZ0h
nGVpKYZsWzt4C9k+9f+3BYM1xWzHkOxE1XBSguSBJ0Z5pUUdHNl/PaDB0W2Q6F6qH2+5AXqJd8Jf
WEUcqR6AJRmsK7T7nH4tS1rlvfmLnR1B9CBaRhPrYz28BBf2H8Esfu5nrhK+oz9XjooMlh3Xwcgm
WIReLmlgWfYlPP199Dd6JKcp+rJ04+EfudvwNk+S09xdkOdc16XXwY3d3kB4ooTvmqH8h+aMaa9p
Wb2RtWy49fUPXiGhV2R9rmWVQ8YuBTgQumwNGjq85hYMLA7EHiCM8mjACGRAWSeXC4zxC2kJB0If
rq79qp8yhMWq76mrKz4wZuY6ka17Oh5ieV0p6qSvgu7/ORboeigoxHQZJHUexdGFsDYpcr3nm2Te
BdbGhb+AMbN9MIMwA0llB+3t3GKvLYB3K/+YdZW/3yvfFZfgJaqFTDyHfuThO62L53bCwIyX7RcH
mmrMisIDlKTbzQEf0/1MMpHMk4m6LB+/6I8S8phcF/InF+ZPFtmq35jD21GW9xXuME+JL5TPeowv
Q0rjWPH54o3MdVXBxxo7Srx6zeKmdJRS7SORiK85YkC5xvQdPBD/5610PTjiNX3b4PvyDDU6/J/O
cNIjiPmjjvJp3cBZlSRLDYGd7M4uD35RQCBGEGqoIjTT/rrZgtTvdJWZ2dCPf+bw8WWT8R0emaxW
1nqzRioztc0KpWUtGUjHtaeL1xrU6DTGH02gf7V3kNBxwZtDZg3Nba/2ddhiMm0behWpG0wKJytw
l97ehGaGdG7hhMscQUcqndlrshkXVIgBHWZo5ktA6CgNsVhWX0eNE1blTr4iKf85ISpo4/iPuvRh
kowxYSMLUZ+kWdGEDtN+pY5Z04JFe2lzIiiYTtne52ooMLEZfAeiBvvAeiAuJHzNFrjdLqZBsG4T
/A3+xG0nteJJlivLWQFIZ1j53gjNAbvUfQcDgUe3hbt/xRCFqvhiAx16CG9QaGS5BgdS5JcEymDw
e0G5U4q/Pk5CIZevd9QR61BilAZm2N+seegtUydyNPNxvgI58xhIQLfNr6VyPZigOeY2MndZXOBf
4ArLeFAxC4xM+ZCJdvMxwpaeXuLb+qKGHfPIfGh0rnyXV7rl2XCPfMVt6fnhWsmXfc1IUnbzLdKH
KvP+2mR7Wf+4YRM6xn586sZpQLMeg+L88aO+7GGJb5LWt5SXhRjWoa3pg9quYu9res8GasNo5Kwu
kXW87Z7z/Text06XKvGfoiRklscVa09UWDOPODJqSUytE5LmdKhesSG5PiHTjUZfhpuzBpasHoH9
5euy1/dCQF15u/AhLk0BMRhoFyAC6o/9dQcJzsRfVoEGSIVlLVxnUBEKWMF/KccaQTQ4BAqT6fxp
CdmZC2R4V8LuG0eho/htzNBAhGcMf/NKVjwsAZoHLq73jqeoq3A2Xac3OeYAGBtTt3OGjVXj7xwz
8CQ5T9lvVqsDbB4tPOphRlYg+wBYL08MkeBuS5scmfFxS5SmFSZLjAVej+fMiMrdnAQqOd9iDffe
bzLHpdBjHgnhSmGypaeNIymUxs5v4Y60d1Nnqp8A+/RLro0unCLhjM8Lv7A3/7BMczM8SgiVV5zM
vFCM6QjgRtK1y1eOU46aCiFCMD16a3nO+xevVsQK1Zca83d3s21N6q4KA93AAcGAZh82BHVuccTq
cRoNTRUhjoNuHvgwT4X7HIHZzrQJW6ssnZgHp/Wz8T4dIQ5bH0Jpt5vj9HVXqnq+uAG631KsEOBZ
n5ROfJf3b/F8XKFjfaqP1zL3gfmcY+2q9KpJCX/2GM2e3wNi0p0mKzVhu8TKHV2MsnEf+eKBl4hN
0+CnpDCfsF4v1O3hzg7oFJcaTs4YMyqqeUe30SH/WfrRQ1Hlt6rxvU5LQGt9xSTeX0Xsx2LTwTbi
g9LT1rC68vqXgoMlraNus3cbNVykbATrOnVhG11AcpLhR5D0Xfng+jV0pZ9QuehFXyCrQlGozLFf
OAEnFodN2ZVPlROZTH/mohcewdURv9WsOO/tZHS6pieChfHRjRLaYmUbuKSVzCPFcp0UY7vKCVKw
arKe/1SYZw1YeMtl2sxkYTlkHlklPw7r16UANAjEBAorY9gyFCdDCmXw+pXFEVzkiIUDn8Vmjz8/
trGOWZzXW3V3+ZDbD+dpITKRnK9R82Q35gsUs7vtP/5nPoPF7jFUtLZWpuZcbsKGttae+cyBdKci
vjhjnbNPY0/IfXKkacDa85zG8o2kLPVxcbqbH3cUxpefWddXAZ1nVxl8CQ4M5x1WPTTp1VB31FPj
oeXjUe+RoWLJjQLC9OwZe9wk39zsnWid4o/tje0JNkr5/Rukc1Gxb1QTTJYc+kawiZU+oPyeaK3B
6v0Hm4CQUwmQSmYkmtr27940+TnoV9+MrWTe+LK2rY3QnatF7RFy4LYMuuU/Qy02FJS/ljFgLjeB
Z/mH9/EZTdkTn2kWEVucw+ClVvDzunANFwrICN1F6alpKumAsMG1TB3gizO9G1GVCUki2gK+fmbb
P4MJb4FhW+8lpoKP/lki2+o9L+gjCd2EEWHRc+eubR9woW8zDU5lDZpTmemdtkW6/K2XgGFXOWRL
5nbwuzhiQcZ5SwzW4vjWviPcEXsTTVeRG2083XD0n4/w2r28JqyE6RsbToukVWENW5ymscZjnckq
8WSFynLq9yIVaQDGx7ItzXnML46yHtM44XVK0npzavsioOLhxZhttTn0VS/gT6jiJeH+dHBufwYh
QNN8sEauGHKpHPaW2kCUPPL6yrWRl9yQRbmre5MIdxlYVH0BOrb+cvs5VxFxvwx0RzqPPKCgw3q4
SNZPer8zXLPtId87gAQumnuMhxsPEqjcTNw+kv48oJ0L/o1d/eMqWEREehC0O2RJshg4HBxwVKE1
r8qXhEcaIpUaUhdG9Zb99JNMOymdTkTKfWHmV5j3GThlguuwpGeiAzJ1076kYFeQ79Xa+yNxVZJq
cuSTyjgNI1cfrmfiHxLPX9pf2JJ27hz6Hl3K3dCde7xLMq37CDVIS+1kCKrQ0riKwnIKH3hSVMc0
ZMBLq0aW2yvITCo1/KNovM7SOBQTzKT+M2WUBydbdQj4s7Tt4LA7wWCKHkQ+Y7cDVnD5lvWPEGhN
F2VjlKiJgYlR4WkNlHQi/aJg0L9TsDlb6box+uYvvxYepG/Oj9aPuXF8RvpoL3FgsovCt8pPjP3n
0340TrjvI/1fGPiMQG6j0bB7LLvDEQyz8Yk2S4V7AT6sa7/LNsF3s0XUHVoUfQp6lTDmdfmSJaxI
XxWfJRnknkvbwLYhBDkvyfX9pn+Mm4RMeoCW5tE4nm2gevFL+iepYDphBlup3gw2efBL6dnx7V7H
M6KaD0Vf9VtJGMdr8jcWn1QqzyMNol/i0RH+KnQGpoi+C5xtJSEtwAkDYF4TlpRfJXmeaylsd9Mw
KyRnzhmJViflJHsBdz1VmHlHPasJLyI0R88iS9ICX0JzmS/xZ3Ow3w7xNaGgIfg3AbgMOOqJCRr3
4Tq/KpN3bfvKDsDxEHwDMKxEhR5HVDb59bR/1WYKh9S2YLIoInU0LPXpqhVB7nQYNOBc4Z5iNZVq
WFhOQfYlcPwQmpa/H31rjT26kx2a4K9bIBLj2hsDQ8z5/TyIOJwbPg6kRR0wzi8O9C6OEFLDWlv0
14Xq+7grjVic+vth0uzO/mtelQPfdNWQNDbmvPrziJGLbKufTsqpK/L7o5EsNubgv6N25HSO8Xzc
Yq7u9ZPa0+vRnJhWQ/eHPiH1TM1OYBBVhulFGFJChsCJx+Fxw0rf/1vq2646rxidQkmU6FeJsY0c
2s70Ca6nZvXV2E2sfebxzzTkps2WLewUzj2lx/3WipIZtVBL5hJVQa1K+qPG984ifySzvPuhzB04
Or6f2xJMX5cNZn/Fr9MfgE/VbiYdwtB9/BwKJoFjR0z0Y7I2YZ1yBBLLmSazZS2gcDJWsXCK+B4O
adaDvWjj3ny+pkaFdUQzIfCYQefYdBH3xMq9GVjqNR0cnH0vgZgz1KTZuoiWL5KJXnYD/ihJ1Afw
mOQ4yMbzaX18c7pt+7WlcLniTh9UG3dTVm1dsXgVONt37XRdZIgK3gPU+itJDwDiBJCy3pRtsnYz
RHpCcJ93TaOWDM/OUybjN6yBBbMY+WES6UPZcOOmd8LkxppgVrlj30bJjDIe96rpLoXhD3Di72wJ
Poyt1GxBrQSRAfQ5+LhmDUbefgbwGzOopou8i5oVbk0xUARthYflJHfkLdPt9yrvH57DFML4oaeI
ehw176xA7k9IE0PPwf/dBbg7DCd5TPVLwrWmzp11WCRNdZEWhRigFZF3rI1eHyp0s5xHdJ5CDJ/H
/JDGxmu+JfEEqSRxXG+qc0QdJMKaBcsdfSClctn/O+cFWDiGwiYD6BsT/bbhVOO10v9M+8IJDpUn
bppLyvg7bWoDJxSMEtojD72RmaFkadkxMxq7avOwRiURzNcLFw7MicKPg3OrG98fM4UdMhQIQP/8
Cllx3GDKnIdQaw==
`protect end_protected
